
module routing_engine_CLOCKED ( port_dest, clk, rst, control, done );
  input [31:0] port_dest;
  output [19:0] control;
  input clk, rst;
  output done;
  wire   \dst[0][2] , \dst[0][1] , \dst[0][0] , \dst[1][2] , \dst[1][1] ,
         \dst[1][0] , \dst[2][2] , \dst[2][1] , \dst[2][0] , \dst[3][2] ,
         \dst[3][0] , \dst[4][2] , \dst[4][1] , \dst[4][0] , \dst[5][2] ,
         \dst[5][1] , \dst[5][0] , \dst[6][2] , \dst[6][1] , \dst[6][0] ,
         \dst[7][1] , \dst[7][0] , \stage_1_output[0][1] ,
         \stage_1_output[0][2] , \stage_1_output[1][2] ,
         \stage_1_output[2][1] , \stage_1_output[2][2] ,
         \stage_1_output[3][2] , \stage_1_output[4][1] , N1614, N1615, N1616,
         N1618, n1, n2, n5, n8, n11, n13, n276, n277, n386, n388, n391, n397,
         n398, n400, n401, n403, n752, n754, n756, n757, n758, n765, n766,
         n785, n799, \control[19] , n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n3, n4, n6, n7, n9, n10, n12, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343;
  assign control[13] = \control[19] ;
  assign control[15] = \control[19] ;
  assign control[19] = \control[19] ;

  DFD1 \stage_1_output_reg[6][1]  ( .D(N1618), .CP(clk), .QN(n343) );
  EDFQD1 \dst_reg[2][0]  ( .D(n2), .E(n785), .CP(clk), .Q(\dst[2][0] ) );
  EDFQD1 \dst_reg[4][0]  ( .D(n1), .E(n1117), .CP(clk), .Q(\dst[4][0] ) );
  EDFQD1 \dst_reg[4][2]  ( .D(n276), .E(n1117), .CP(clk), .Q(\dst[4][2] ) );
  EDFQD1 \dst_reg[2][2]  ( .D(n799), .E(n785), .CP(clk), .Q(\dst[2][2] ) );
  EDFQD1 \dst_reg[2][1]  ( .D(n1118), .E(n785), .CP(clk), .Q(\dst[2][1] ) );
  DFKCNQD1 \stage_1_output_reg[4][1]  ( .CN(done), .D(n401), .CP(clk), .Q(
        \stage_1_output[4][1] ) );
  DFQD1 \dst_reg[0][1]  ( .D(n758), .CP(clk), .Q(\dst[0][1] ) );
  DFQD1 \dst_reg[5][1]  ( .D(n1115), .CP(clk), .Q(\dst[5][1] ) );
  DFQD1 \dst_reg[5][0]  ( .D(n391), .CP(clk), .Q(\dst[5][0] ) );
  DFQD1 \dst_reg[6][1]  ( .D(n766), .CP(clk), .Q(\dst[6][1] ) );
  DFQD1 \dst_reg[1][2]  ( .D(n1113), .CP(clk), .Q(\dst[1][2] ) );
  DFQD1 \dst_reg[0][2]  ( .D(n757), .CP(clk), .Q(\dst[0][2] ) );
  DFQD1 \dst_reg[7][0]  ( .D(n386), .CP(clk), .Q(\dst[7][0] ) );
  DFQD1 \dst_reg[3][2]  ( .D(n13), .CP(clk), .Q(\dst[3][2] ) );
  DFQD1 \dst_reg[0][0]  ( .D(n403), .CP(clk), .Q(\dst[0][0] ) );
  DFQD1 \dst_reg[1][1]  ( .D(n401), .CP(clk), .Q(\dst[1][1] ) );
  DFQD1 \dst_reg[1][0]  ( .D(n400), .CP(clk), .Q(\dst[1][0] ) );
  DFQD1 \dst_reg[3][0]  ( .D(n397), .CP(clk), .Q(\dst[3][0] ) );
  DFQD1 \dst_reg[6][0]  ( .D(n388), .CP(clk), .Q(\dst[6][0] ) );
  DFQD1 \dst_reg[5][2]  ( .D(n1114), .CP(clk), .Q(\dst[5][2] ) );
  DFQD1 \dst_reg[7][1]  ( .D(n1116), .CP(clk), .Q(\dst[7][1] ) );
  DFXQD1 \stage_1_output_reg[0][2]  ( .DB(n400), .DA(n403), .SA(done), .CP(clk), .Q(\stage_1_output[0][2] ) );
  DFXQD1 \stage_1_output_reg[1][2]  ( .DB(n397), .DA(n398), .SA(n1112), .CP(
        clk), .Q(\stage_1_output[1][2] ) );
  DFQD1 \stage_1_output_reg[0][1]  ( .D(n758), .CP(clk), .Q(
        \stage_1_output[0][1] ) );
  DFQD1 \stage_1_output_reg[2][1]  ( .D(N1615), .CP(clk), .Q(
        \stage_1_output[2][1] ) );
  DFQD1 \dst_reg[6][2]  ( .D(n765), .CP(clk), .Q(\dst[6][2] ) );
  DFQD1 \stage_1_output_reg[2][2]  ( .D(N1614), .CP(clk), .Q(
        \stage_1_output[2][2] ) );
  DFQD1 \stage_1_output_reg[3][2]  ( .D(N1616), .CP(clk), .Q(
        \stage_1_output[3][2] ) );
  EDFQD1 \dst_reg[4][1]  ( .D(n277), .E(n1117), .CP(clk), .Q(\dst[4][1] ) );
  DFQD1 \stage_0_sw_ctl_reg[1]  ( .D(n756), .CP(clk), .Q(control[18]) );
  DFQD1 \stage_0_sw_ctl_reg[2]  ( .D(n754), .CP(clk), .Q(control[17]) );
  DFQD1 \stage_1_sw_ctl_reg[3]  ( .D(n5), .CP(clk), .Q(control[12]) );
  DFQD1 \stage_1_sw_ctl_reg[1]  ( .D(n752), .CP(clk), .Q(control[14]) );
  DFQD1 \stage_0_sw_ctl_reg[3]  ( .D(n8), .CP(clk), .Q(control[16]) );
  DFKCNQD1 \stage_1_output_reg[4][0]  ( .CN(done), .D(n1113), .CP(clk), .Q(
        control[9]) );
  DFQD1 \stage_1_output_reg[0][0]  ( .D(n757), .CP(clk), .Q(control[11]) );
  DFXQD1 \stage_1_output_reg[5][0]  ( .DB(n11), .DA(n13), .SA(n1112), .CP(clk), 
        .Q(control[8]) );
  DFXQD1 \stage_1_output_reg[1][0]  ( .DB(n13), .DA(n11), .SA(n1112), .CP(clk), 
        .Q(control[10]) );
  MUX2ND1 U422 ( .I0(n66), .I1(n67), .S(control[7]), .ZN(control[3]) );
  MUX2ND1 U423 ( .I0(n68), .I1(n69), .S(control[6]), .ZN(control[1]) );
  MUX2ND1 U424 ( .I0(n69), .I1(n68), .S(control[6]), .ZN(control[0]) );
  CKMUX2D1 U425 ( .I0(\stage_1_output[2][1] ), .I1(\stage_1_output[0][1] ), 
        .S(control[11]), .Z(control[6]) );
  MUX2ND1 U426 ( .I0(n67), .I1(n66), .S(control[7]), .ZN(control[2]) );
  MUX2ND1 U427 ( .I0(n343), .I1(n65), .S(control[9]), .ZN(control[4]) );
  CKMUX2D1 U428 ( .I0(\stage_1_output[0][1] ), .I1(\stage_1_output[2][1] ), 
        .S(control[11]), .Z(control[7]) );
  MUX2ND1 U429 ( .I0(n65), .I1(n343), .S(control[9]), .ZN(control[5]) );
  TIEH U430 ( .Z(done) );
  TIEL U431 ( .ZN(\control[19] ) );
  CKND0 U432 ( .I(n3), .ZN(n799) );
  CKND0 U433 ( .I(n1112), .ZN(n756) );
  CKND0 U434 ( .I(n4), .ZN(n5) );
  MUX3D0 U435 ( .I0(port_dest[28]), .I1(n6), .I2(\dst[0][0] ), .S0(n7), .S1(n9), .Z(n403) );
  INR4D0 U436 ( .A1(n10), .B1(n12), .B2(n14), .B3(n15), .ZN(n6) );
  NR2D0 U437 ( .A1(n16), .A2(n17), .ZN(n15) );
  MUX3D0 U438 ( .I0(port_dest[25]), .I1(n18), .I2(\dst[1][1] ), .S0(n19), .S1(
        n20), .Z(n401) );
  OAI211D0 U439 ( .A1(n21), .A2(n22), .B(n23), .C(n24), .ZN(n18) );
  CKND0 U440 ( .I(n25), .ZN(n23) );
  MUX3D0 U441 ( .I0(port_dest[24]), .I1(n26), .I2(\dst[1][0] ), .S0(n19), .S1(
        n20), .Z(n400) );
  CKND0 U442 ( .I(n27), .ZN(n20) );
  NR3D0 U443 ( .A1(n28), .A2(n29), .A3(n25), .ZN(n26) );
  MUX2D0 U444 ( .I0(\dst[2][0] ), .I1(n2), .S(n785), .Z(n398) );
  MUX3D0 U445 ( .I0(port_dest[16]), .I1(n30), .I2(\dst[3][0] ), .S0(n31), .S1(
        n32), .Z(n397) );
  AOI211D0 U446 ( .A1(n33), .A2(n34), .B(n35), .C(n36), .ZN(n30) );
  CKND0 U447 ( .I(n37), .ZN(n36) );
  CKND0 U448 ( .I(n38), .ZN(n391) );
  MUX2D0 U449 ( .I0(n39), .I1(port_dest[20]), .S(port_dest[23]), .Z(n2) );
  AOI211D0 U450 ( .A1(n40), .A2(n41), .B(n42), .C(n43), .ZN(n39) );
  CKND0 U451 ( .I(n44), .ZN(n42) );
  AO221D0 U452 ( .A1(n45), .A2(n31), .B1(\dst[3][2] ), .B2(n32), .C(n46), .Z(
        n13) );
  AN3D0 U453 ( .A1(n47), .A2(n48), .A3(n49), .Z(n32) );
  CKND2D0 U454 ( .A1(n49), .A2(n48), .ZN(n45) );
  CKND2D0 U455 ( .A1(n50), .A2(n51), .ZN(n48) );
  IAO21D0 U456 ( .A1(n52), .A2(n53), .B(n35), .ZN(n49) );
  OAI22D0 U457 ( .A1(n52), .A2(n54), .B1(n55), .B2(n56), .ZN(n35) );
  CKND0 U458 ( .I(n51), .ZN(n55) );
  CKND0 U459 ( .I(n57), .ZN(n1114) );
  OAI221D0 U460 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .C(n62), .ZN(n1112)
         );
  AN2D0 U461 ( .A1(n63), .A2(n64), .Z(n62) );
  CKND0 U462 ( .I(\stage_1_output[4][1] ), .ZN(n65) );
  MUX2ND0 U463 ( .I0(\stage_1_output[0][2] ), .I1(\stage_1_output[2][2] ), .S(
        control[11]), .ZN(n66) );
  MUX2ND0 U464 ( .I0(\stage_1_output[1][2] ), .I1(\stage_1_output[3][2] ), .S(
        control[10]), .ZN(n67) );
  MUX2ND0 U465 ( .I0(\stage_1_output[2][2] ), .I1(\stage_1_output[0][2] ), .S(
        control[11]), .ZN(n68) );
  MUX2ND0 U466 ( .I0(\stage_1_output[3][2] ), .I1(\stage_1_output[1][2] ), .S(
        control[10]), .ZN(n69) );
  MUX3ND0 U467 ( .I0(n70), .I1(n71), .I2(n72), .S0(n8), .S1(n4), .ZN(N1618) );
  CKXOR2D0 U468 ( .A1(n73), .A2(n1113), .Z(n4) );
  OA32D0 U469 ( .A1(n74), .A2(n75), .A3(n76), .B1(\dst[1][2] ), .B2(n27), .Z(
        n1113) );
  ND4D0 U470 ( .A1(n77), .A2(n78), .A3(n79), .A4(n22), .ZN(n27) );
  NR2D0 U471 ( .A1(n80), .A2(n25), .ZN(n79) );
  NR2D0 U472 ( .A1(n81), .A2(n21), .ZN(n25) );
  NR2D0 U473 ( .A1(port_dest[27]), .A2(n77), .ZN(n74) );
  AOI21D0 U474 ( .A1(n82), .A2(n83), .B(n28), .ZN(n77) );
  MOAI22D0 U475 ( .A1(n24), .A2(n84), .B1(n82), .B2(n85), .ZN(n28) );
  CKND0 U476 ( .I(n86), .ZN(n82) );
  MUX2ND0 U477 ( .I0(n57), .I1(n87), .S(n754), .ZN(n73) );
  MUX2ND0 U478 ( .I0(n1115), .I1(n88), .S(n754), .ZN(n72) );
  CKND0 U479 ( .I(n89), .ZN(n1115) );
  MUX2ND0 U480 ( .I0(n90), .I1(n91), .S(n752), .ZN(N1616) );
  MUX3ND0 U481 ( .I0(n92), .I1(n89), .I2(n93), .S0(n754), .S1(n752), .ZN(N1615) );
  MUX2ND0 U482 ( .I0(n766), .I1(n1116), .S(n8), .ZN(n93) );
  CKND0 U483 ( .I(n70), .ZN(n1116) );
  MUX2ND0 U484 ( .I0(n94), .I1(\dst[7][1] ), .S(n95), .ZN(n70) );
  CKND2D0 U485 ( .A1(n96), .A2(n97), .ZN(n94) );
  OAI21D0 U486 ( .A1(n98), .A2(n99), .B(n100), .ZN(n97) );
  CKND0 U487 ( .I(n101), .ZN(n99) );
  CKND0 U488 ( .I(n71), .ZN(n766) );
  AOI211D0 U489 ( .A1(\dst[5][1] ), .A2(n102), .B(n103), .C(n104), .ZN(n89) );
  AOI31D0 U490 ( .A1(n105), .A2(n106), .A3(n107), .B(n108), .ZN(n104) );
  MUX2ND0 U491 ( .I0(n91), .I1(n90), .S(n752), .ZN(N1614) );
  XNR2D0 U492 ( .A1(n109), .A2(n757), .ZN(n752) );
  MUX2ND0 U493 ( .I0(n87), .I1(n57), .S(n754), .ZN(n109) );
  AOI221D0 U494 ( .A1(n110), .A2(n111), .B1(\dst[5][2] ), .B2(n102), .C(n112), 
        .ZN(n57) );
  IND2D0 U495 ( .A1(n113), .B1(n114), .ZN(n111) );
  MUX2ND0 U496 ( .I0(n388), .I1(n386), .S(n8), .ZN(n90) );
  OAI21D0 U497 ( .A1(n115), .A2(n116), .B(n117), .ZN(n8) );
  MUX4ND0 U498 ( .I0(n118), .I1(n119), .I2(n120), .I3(n121), .S0(n122), .S1(
        n71), .ZN(n117) );
  IAO21D0 U499 ( .A1(\dst[6][2] ), .A2(n123), .B(n124), .ZN(n122) );
  AOI211D0 U500 ( .A1(n125), .A2(n126), .B(n127), .C(n128), .ZN(n124) );
  CKND2D0 U501 ( .A1(n63), .A2(n129), .ZN(n121) );
  IND2D0 U502 ( .A1(n130), .B1(n60), .ZN(n120) );
  CKND2D0 U503 ( .A1(n64), .A2(n131), .ZN(n119) );
  CKND2D0 U504 ( .A1(n58), .A2(n132), .ZN(n118) );
  XNR2D0 U505 ( .A1(n765), .A2(n133), .ZN(n116) );
  OA32D0 U506 ( .A1(n134), .A2(n127), .A3(n128), .B1(\dst[6][2] ), .B2(n123), 
        .Z(n765) );
  NR2D0 U507 ( .A1(n135), .A2(port_dest[7]), .ZN(n134) );
  XNR2D0 U508 ( .A1(n71), .A2(n758), .ZN(n115) );
  OAI22D0 U509 ( .A1(\dst[6][1] ), .A2(n123), .B1(n128), .B2(n136), .ZN(n71)
         );
  MUX2ND0 U510 ( .I0(n137), .I1(n138), .S(n125), .ZN(n136) );
  NR2D0 U511 ( .A1(n139), .A2(n140), .ZN(n138) );
  IAO21D0 U512 ( .A1(n141), .A2(n142), .B(n143), .ZN(n140) );
  CKND0 U513 ( .I(n144), .ZN(n123) );
  AO21D0 U514 ( .A1(\dst[7][0] ), .A2(n95), .B(n145), .Z(n386) );
  MUX2ND0 U515 ( .I0(n146), .I1(n147), .S(n100), .ZN(n145) );
  NR2D0 U516 ( .A1(n148), .A2(n149), .ZN(n147) );
  NR4D0 U517 ( .A1(n98), .A2(n150), .A3(n151), .A4(n152), .ZN(n148) );
  AN4D0 U518 ( .A1(n153), .A2(n154), .A3(n101), .A4(n155), .Z(n95) );
  INR4D0 U519 ( .A1(n156), .B1(port_dest[3]), .B2(n149), .B3(n151), .ZN(n155)
         );
  INR2D0 U520 ( .A1(n157), .B1(n158), .ZN(n151) );
  CKND0 U521 ( .I(n159), .ZN(n149) );
  IND4D0 U522 ( .A1(n128), .B1(n98), .B2(n160), .B3(n154), .ZN(n159) );
  AN3D0 U523 ( .A1(n158), .A2(n156), .A3(n157), .Z(n98) );
  AOI21D0 U524 ( .A1(n161), .A2(n141), .B(n162), .ZN(n157) );
  OAI21D0 U525 ( .A1(n141), .A2(n161), .B(n163), .ZN(n158) );
  NR3D0 U526 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n128) );
  CKND2D0 U527 ( .A1(n165), .A2(n166), .ZN(n156) );
  AOI31D0 U528 ( .A1(n167), .A2(n161), .A3(n141), .B(n152), .ZN(n101) );
  OA211D0 U529 ( .A1(port_dest[7]), .A2(n143), .B(n142), .C(n153), .Z(n152) );
  CKND0 U530 ( .I(n162), .ZN(n167) );
  OAI21D0 U531 ( .A1(n168), .A2(n169), .B(n153), .ZN(n162) );
  NR2D0 U532 ( .A1(port_dest[7]), .A2(n143), .ZN(n168) );
  OAI21D0 U533 ( .A1(n165), .A2(n166), .B(n164), .ZN(n154) );
  CKND2D0 U534 ( .A1(n170), .A2(n125), .ZN(n166) );
  INR2D0 U535 ( .A1(n171), .B1(n150), .ZN(n153) );
  NR2D0 U536 ( .A1(n172), .A2(n125), .ZN(n150) );
  OAI21D0 U537 ( .A1(port_dest[7]), .A2(n173), .B(n174), .ZN(n171) );
  MUX3D0 U538 ( .I0(n175), .I1(port_dest[4]), .I2(\dst[6][0] ), .S0(
        port_dest[7]), .S1(n144), .Z(n388) );
  NR4D0 U539 ( .A1(n161), .A2(n126), .A3(n141), .A4(n160), .ZN(n144) );
  AOI31D0 U540 ( .A1(n176), .A2(n177), .A3(n178), .B(n179), .ZN(n160) );
  CKND0 U541 ( .I(n135), .ZN(n126) );
  AOI211D0 U542 ( .A1(n170), .A2(n165), .B(n180), .C(n139), .ZN(n135) );
  OR3D0 U543 ( .A1(n143), .A2(n142), .A3(port_dest[7]), .Z(n161) );
  NR4D0 U544 ( .A1(n173), .A2(n139), .A3(n180), .A4(n181), .ZN(n175) );
  NR2D0 U545 ( .A1(n143), .A2(n169), .ZN(n181) );
  CKND0 U546 ( .I(n142), .ZN(n169) );
  AN2D0 U547 ( .A1(n163), .A2(n182), .Z(n180) );
  CKND0 U548 ( .I(n183), .ZN(n139) );
  IND3D0 U549 ( .A1(n165), .B1(n164), .B2(n170), .ZN(n183) );
  INR2D0 U550 ( .A1(n182), .B1(n163), .ZN(n170) );
  OA21D0 U551 ( .A1(port_dest[11]), .A2(n184), .B(n185), .Z(n163) );
  NR3D0 U552 ( .A1(n141), .A2(n142), .A3(n143), .ZN(n182) );
  OR2D0 U553 ( .A1(n174), .A2(n173), .Z(n143) );
  OA21D0 U554 ( .A1(port_dest[11]), .A2(n186), .B(n187), .Z(n174) );
  AOI21D0 U555 ( .A1(n177), .A2(n188), .B(n189), .ZN(n142) );
  AOI31D0 U556 ( .A1(n188), .A2(n177), .A3(n189), .B(n190), .ZN(n141) );
  AOI21D0 U557 ( .A1(n177), .A2(n176), .B(n178), .ZN(n164) );
  CKND0 U558 ( .I(n191), .ZN(n178) );
  AOI21D0 U559 ( .A1(n177), .A2(n113), .B(n192), .ZN(n165) );
  CKND0 U560 ( .I(n172), .ZN(n173) );
  CKND2D0 U561 ( .A1(n186), .A2(port_dest[11]), .ZN(n172) );
  MUX2D0 U562 ( .I0(n193), .I1(n38), .S(n754), .Z(n91) );
  AN3D0 U563 ( .A1(n131), .A2(n129), .A3(n194), .Z(n754) );
  AOI33D0 U564 ( .A1(n195), .A2(n196), .A3(n58), .B1(n197), .B2(n130), .B3(n60), .ZN(n194) );
  AOI22D0 U565 ( .A1(n3), .A2(n198), .B1(n199), .B2(n200), .ZN(n60) );
  OAI22D0 U566 ( .A1(n277), .A2(n276), .B1(\dst[4][1] ), .B2(n201), .ZN(n130)
         );
  CKND0 U567 ( .I(n61), .ZN(n197) );
  NR2D0 U568 ( .A1(n757), .A2(n758), .ZN(n61) );
  AOI32D0 U569 ( .A1(\dst[2][1] ), .A2(n199), .A3(n202), .B1(n3), .B2(n1118), 
        .ZN(n58) );
  CKND0 U570 ( .I(n132), .ZN(n196) );
  AOI22D0 U571 ( .A1(n203), .A2(\dst[4][1] ), .B1(n204), .B2(n277), .ZN(n132)
         );
  CKND0 U572 ( .I(n59), .ZN(n195) );
  NR2D0 U573 ( .A1(n205), .A2(n757), .ZN(n59) );
  OAI211D0 U574 ( .A1(n758), .A2(n133), .B(n206), .C(n63), .ZN(n129) );
  OAI21D0 U575 ( .A1(n758), .A2(n133), .B(n207), .ZN(n63) );
  MOAI22D0 U576 ( .A1(n1118), .A2(n3), .B1(n200), .B2(\dst[2][2] ), .ZN(n207)
         );
  OAI32D0 U577 ( .A1(n208), .A2(\dst[4][1] ), .A3(n1117), .B1(n277), .B2(n204), 
        .ZN(n206) );
  CKND0 U578 ( .I(\dst[4][2] ), .ZN(n208) );
  IND4D0 U579 ( .A1(n87), .B1(n88), .B2(n209), .B3(n64), .ZN(n131) );
  OAI211D0 U580 ( .A1(n133), .A2(n205), .B(n11), .C(n210), .ZN(n64) );
  NR2D0 U581 ( .A1(n200), .A2(n198), .ZN(n210) );
  CKND0 U582 ( .I(n1118), .ZN(n198) );
  OAI221D0 U583 ( .A1(n211), .A2(n212), .B1(n213), .B2(n214), .C(n215), .ZN(
        n1118) );
  NR2D0 U584 ( .A1(n785), .A2(\dst[2][1] ), .ZN(n200) );
  MUX2ND0 U585 ( .I0(n3), .I1(n199), .S(n202), .ZN(n11) );
  CKND0 U586 ( .I(n785), .ZN(n202) );
  ND4D0 U587 ( .A1(n216), .A2(n217), .A3(n218), .A4(n44), .ZN(n785) );
  CKND2D0 U588 ( .A1(n219), .A2(n220), .ZN(n44) );
  IOA21D0 U589 ( .A1(n218), .A2(n221), .B(n222), .ZN(n220) );
  CKND0 U590 ( .I(\dst[2][2] ), .ZN(n199) );
  NR2D0 U591 ( .A1(n216), .A2(n223), .ZN(n3) );
  CKND2D0 U592 ( .A1(n758), .A2(n757), .ZN(n209) );
  CKND0 U593 ( .I(n133), .ZN(n757) );
  INR3D0 U594 ( .A1(n224), .B1(n225), .B2(n226), .ZN(n133) );
  AOI22D0 U595 ( .A1(n7), .A2(n227), .B1(\dst[0][2] ), .B2(n9), .ZN(n224) );
  CKND0 U596 ( .I(n205), .ZN(n758) );
  AOI211D0 U597 ( .A1(\dst[0][1] ), .A2(n9), .B(n225), .C(n228), .ZN(n205) );
  MUX2ND0 U598 ( .I0(n229), .I1(n230), .S(n7), .ZN(n228) );
  NR2D0 U599 ( .A1(n12), .A2(n231), .ZN(n230) );
  NR2D0 U600 ( .A1(n232), .A2(n9), .ZN(n225) );
  INR4D0 U601 ( .A1(n233), .B1(n234), .B2(n227), .B3(n231), .ZN(n9) );
  NR2D0 U602 ( .A1(n235), .A2(n236), .ZN(n231) );
  OAI21D0 U603 ( .A1(n237), .A2(n16), .B(n10), .ZN(n227) );
  ND3D0 U604 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n10) );
  AN2D0 U605 ( .A1(n17), .A2(n240), .Z(n237) );
  NR2D0 U606 ( .A1(n12), .A2(n241), .ZN(n233) );
  INR3D0 U607 ( .A1(n242), .B1(n14), .B2(n243), .ZN(n12) );
  CKND0 U608 ( .I(n244), .ZN(n14) );
  CKND0 U609 ( .I(n92), .ZN(n88) );
  OAI21D0 U610 ( .A1(\dst[4][1] ), .A2(n1117), .B(n277), .ZN(n92) );
  CKND2D0 U611 ( .A1(n245), .A2(n246), .ZN(n277) );
  MUX2ND0 U612 ( .I0(port_dest[13]), .I1(n247), .S(n248), .ZN(n245) );
  OAI211D0 U613 ( .A1(n249), .A2(n250), .B(n251), .C(n252), .ZN(n247) );
  CKND2D0 U614 ( .A1(n276), .A2(n201), .ZN(n87) );
  CKND0 U615 ( .I(n203), .ZN(n201) );
  NR2D0 U616 ( .A1(n1117), .A2(\dst[4][2] ), .ZN(n203) );
  CKND0 U617 ( .I(n204), .ZN(n276) );
  NR2D0 U618 ( .A1(n253), .A2(n254), .ZN(n204) );
  AOI221D0 U619 ( .A1(\dst[5][0] ), .A2(n102), .B1(port_dest[8]), .B2(
        port_dest[11]), .C(n255), .ZN(n38) );
  IINR4D0 U620 ( .A1(n114), .A2(n106), .B1(n186), .B2(n108), .ZN(n255) );
  CKND0 U621 ( .I(n110), .ZN(n108) );
  NR2D0 U622 ( .A1(n102), .A2(port_dest[11]), .ZN(n110) );
  AN4D0 U623 ( .A1(n188), .A2(n179), .A3(n114), .A4(n256), .Z(n102) );
  AN4D0 U624 ( .A1(n177), .A2(n106), .A3(n105), .A4(n192), .Z(n256) );
  IND2D0 U625 ( .A1(n190), .B1(n188), .ZN(n105) );
  IND2D0 U626 ( .A1(n189), .B1(n188), .ZN(n106) );
  AOI22D0 U627 ( .A1(n257), .A2(n185), .B1(n176), .B2(n191), .ZN(n114) );
  NR2D0 U628 ( .A1(n258), .A2(n259), .ZN(n191) );
  CKND0 U629 ( .I(n107), .ZN(n176) );
  CKND2D0 U630 ( .A1(n113), .A2(n192), .ZN(n107) );
  IOA21D0 U631 ( .A1(n260), .A2(n253), .B(n261), .ZN(n192) );
  NR2D0 U632 ( .A1(n184), .A2(n185), .ZN(n113) );
  NR2D0 U633 ( .A1(n260), .A2(n253), .ZN(n185) );
  CKND0 U634 ( .I(n184), .ZN(n257) );
  ND3D0 U635 ( .A1(n190), .A2(n189), .A3(n188), .ZN(n184) );
  OAI21D0 U636 ( .A1(port_dest[15]), .A2(n249), .B(n262), .ZN(n189) );
  OAI31D0 U637 ( .A1(n249), .A2(port_dest[15]), .A3(n262), .B(n263), .ZN(n190)
         );
  CKND0 U638 ( .I(n264), .ZN(n249) );
  ND3D0 U639 ( .A1(n265), .A2(n246), .A3(n50), .ZN(n179) );
  CKND2D0 U640 ( .A1(n259), .A2(n258), .ZN(n246) );
  CKND0 U641 ( .I(n266), .ZN(n258) );
  INR2D0 U642 ( .A1(n267), .B1(port_dest[15]), .ZN(n259) );
  NR2D0 U643 ( .A1(n187), .A2(n186), .ZN(n188) );
  AN2D0 U644 ( .A1(n268), .A2(port_dest[15]), .Z(n186) );
  OA21D0 U645 ( .A1(n268), .A2(port_dest[15]), .B(n269), .Z(n187) );
  OAI21D0 U646 ( .A1(\dst[4][0] ), .A2(n1117), .B(n1), .ZN(n193) );
  MUX2D0 U647 ( .I0(n270), .I1(port_dest[12]), .S(port_dest[15]), .Z(n1) );
  INR3D0 U648 ( .A1(n251), .B1(n271), .B2(n268), .ZN(n270) );
  CKND2D0 U649 ( .A1(n262), .A2(n264), .ZN(n251) );
  CKND0 U650 ( .I(n272), .ZN(n262) );
  IIND4D0 U651 ( .A1(n271), .A2(n261), .B1(n253), .B2(n273), .ZN(n1117) );
  CKND2D0 U652 ( .A1(n50), .A2(n265), .ZN(n273) );
  ND3D0 U653 ( .A1(n56), .A2(n31), .A3(n51), .ZN(n265) );
  IAO21D0 U654 ( .A1(n221), .A2(n215), .B(n217), .ZN(n50) );
  IOA21D0 U655 ( .A1(n84), .A2(n76), .B(n80), .ZN(n217) );
  OA21D0 U656 ( .A1(n239), .A2(n232), .B(n241), .Z(n80) );
  AN4D0 U657 ( .A1(n274), .A2(n275), .A3(n278), .A4(n279), .Z(n241) );
  AOI33D0 U658 ( .A1(port_dest[28]), .A2(n226), .A3(port_dest[29]), .B1(
        port_dest[4]), .B2(n127), .B3(port_dest[5]), .ZN(n279) );
  AOI33D0 U659 ( .A1(port_dest[24]), .A2(n75), .A3(port_dest[25]), .B1(
        port_dest[20]), .B2(n223), .B3(port_dest[21]), .ZN(n278) );
  AOI33D0 U660 ( .A1(port_dest[16]), .A2(n46), .A3(port_dest[17]), .B1(
        port_dest[12]), .B2(n254), .B3(port_dest[13]), .ZN(n275) );
  AOI33D0 U661 ( .A1(port_dest[2]), .A2(port_dest[0]), .A3(n280), .B1(
        port_dest[8]), .B2(port_dest[10]), .B3(n103), .ZN(n274) );
  NR2D0 U662 ( .A1(n281), .A2(port_dest[15]), .ZN(n253) );
  OAI21D0 U663 ( .A1(n281), .A2(n260), .B(n252), .ZN(n271) );
  CKND2D0 U664 ( .A1(n266), .A2(n267), .ZN(n252) );
  NR3D0 U665 ( .A1(n261), .A2(n282), .A3(n281), .ZN(n267) );
  AOI21D0 U666 ( .A1(n54), .A2(n47), .B(n53), .ZN(n261) );
  CKND0 U667 ( .I(n283), .ZN(n53) );
  AOI21D0 U668 ( .A1(n31), .A2(n51), .B(n56), .ZN(n266) );
  CKND2D0 U669 ( .A1(n221), .A2(n215), .ZN(n56) );
  ND3D0 U670 ( .A1(n218), .A2(n222), .A3(n216), .ZN(n215) );
  NR2D0 U671 ( .A1(n84), .A2(n76), .ZN(n221) );
  NR2D0 U672 ( .A1(n24), .A2(port_dest[27]), .ZN(n76) );
  OR3D0 U673 ( .A1(n85), .A2(n83), .A3(n86), .Z(n24) );
  CKND2D0 U674 ( .A1(n239), .A2(n232), .ZN(n84) );
  CKND2D0 U675 ( .A1(n284), .A2(n240), .ZN(n232) );
  AN4D0 U676 ( .A1(n285), .A2(n286), .A3(n287), .A4(n288), .Z(n239) );
  AOI33D0 U677 ( .A1(n226), .A2(n289), .A3(port_dest[29]), .B1(n127), .B2(n290), .B3(port_dest[5]), .ZN(n288) );
  AOI33D0 U678 ( .A1(n75), .A2(n291), .A3(port_dest[25]), .B1(n223), .B2(n292), 
        .B3(port_dest[21]), .ZN(n287) );
  AOI33D0 U679 ( .A1(n46), .A2(n293), .A3(port_dest[17]), .B1(n254), .B2(n294), 
        .B3(port_dest[13]), .ZN(n286) );
  AOI33D0 U680 ( .A1(port_dest[2]), .A2(n146), .A3(n280), .B1(port_dest[10]), 
        .B2(n295), .B3(n103), .ZN(n285) );
  NR3D0 U681 ( .A1(n283), .A2(n296), .A3(n52), .ZN(n51) );
  AOI21D0 U682 ( .A1(n222), .A2(n216), .B(n218), .ZN(n283) );
  OAI31D0 U683 ( .A1(n86), .A2(port_dest[27]), .A3(n85), .B(n83), .ZN(n218) );
  NR2D0 U684 ( .A1(n240), .A2(n284), .ZN(n83) );
  INR3D0 U685 ( .A1(n17), .B1(port_dest[31]), .B2(n16), .ZN(n284) );
  CKND0 U686 ( .I(n238), .ZN(n16) );
  ND4D0 U687 ( .A1(n297), .A2(n298), .A3(n299), .A4(n300), .ZN(n240) );
  AOI33D0 U688 ( .A1(n112), .A2(n301), .A3(port_dest[8]), .B1(n226), .B2(n229), 
        .B3(port_dest[28]), .ZN(n300) );
  AOI33D0 U689 ( .A1(n127), .A2(n137), .A3(port_dest[4]), .B1(n75), .B2(n302), 
        .B3(port_dest[24]), .ZN(n299) );
  AOI33D0 U690 ( .A1(n223), .A2(n214), .A3(port_dest[20]), .B1(n46), .B2(n303), 
        .B3(port_dest[16]), .ZN(n298) );
  AOI33D0 U691 ( .A1(n254), .A2(n304), .A3(port_dest[12]), .B1(port_dest[0]), 
        .B2(n305), .B3(port_dest[2]), .ZN(n297) );
  CKND0 U692 ( .I(n282), .ZN(n260) );
  NR2D0 U693 ( .A1(n54), .A2(n47), .ZN(n282) );
  NR2D0 U694 ( .A1(n52), .A2(port_dest[19]), .ZN(n47) );
  ND4D0 U695 ( .A1(n306), .A2(n307), .A3(n34), .A4(n37), .ZN(n52) );
  CKND0 U696 ( .I(n296), .ZN(n54) );
  NR2D0 U697 ( .A1(n222), .A2(n216), .ZN(n296) );
  INR2D0 U698 ( .A1(n219), .B1(port_dest[23]), .ZN(n216) );
  AN2D0 U699 ( .A1(n41), .A2(n211), .Z(n219) );
  NR2D0 U700 ( .A1(n40), .A2(n308), .ZN(n211) );
  OAI21D0 U701 ( .A1(port_dest[27]), .A2(n86), .B(n85), .ZN(n222) );
  AOI21D0 U702 ( .A1(n7), .A2(n238), .B(n17), .ZN(n85) );
  ND4D0 U703 ( .A1(n309), .A2(n310), .A3(n311), .A4(n312), .ZN(n17) );
  AOI33D0 U704 ( .A1(n293), .A2(n303), .A3(n46), .B1(n294), .B2(n304), .B3(
        n254), .ZN(n312) );
  INR2D0 U705 ( .A1(port_dest[14]), .B1(n248), .ZN(n254) );
  AN2D0 U706 ( .A1(port_dest[18]), .A2(port_dest[19]), .Z(n46) );
  AOI33D0 U707 ( .A1(n291), .A2(n302), .A3(n75), .B1(n292), .B2(n214), .B3(
        n223), .ZN(n311) );
  INR2D0 U708 ( .A1(port_dest[22]), .B1(n213), .ZN(n223) );
  AN2D0 U709 ( .A1(port_dest[26]), .A2(port_dest[27]), .Z(n75) );
  AOI33D0 U710 ( .A1(n290), .A2(n137), .A3(n127), .B1(n289), .B2(n229), .B3(
        n226), .ZN(n310) );
  INR2D0 U711 ( .A1(port_dest[30]), .B1(n7), .ZN(n226) );
  AN2D0 U712 ( .A1(port_dest[6]), .A2(port_dest[7]), .Z(n127) );
  AOI33D0 U713 ( .A1(n295), .A2(n301), .A3(n112), .B1(n305), .B2(n146), .B3(
        port_dest[2]), .ZN(n309) );
  NR2D0 U714 ( .A1(n177), .A2(n313), .ZN(n112) );
  NR2D0 U715 ( .A1(n236), .A2(n314), .ZN(n238) );
  ND3D0 U716 ( .A1(n22), .A2(n81), .A3(n315), .ZN(n86) );
  ND3D0 U717 ( .A1(n250), .A2(n272), .A3(n264), .ZN(n281) );
  NR2D0 U718 ( .A1(n269), .A2(n268), .ZN(n264) );
  NR2D0 U719 ( .A1(n37), .A2(n31), .ZN(n268) );
  AOI21D0 U720 ( .A1(n31), .A2(n37), .B(n34), .ZN(n269) );
  CKND2D0 U721 ( .A1(n33), .A2(n316), .ZN(n272) );
  CKND0 U722 ( .I(n263), .ZN(n250) );
  IAO21D0 U723 ( .A1(n33), .A2(n316), .B(n306), .ZN(n263) );
  OAI21D0 U724 ( .A1(n40), .A2(n212), .B(n308), .ZN(n306) );
  AOI21D0 U725 ( .A1(n81), .A2(n78), .B(n22), .ZN(n308) );
  OAI21D0 U726 ( .A1(port_dest[31]), .A2(n236), .B(n314), .ZN(n22) );
  CKND0 U727 ( .I(n235), .ZN(n314) );
  ND4D0 U728 ( .A1(n317), .A2(n318), .A3(n319), .A4(n320), .ZN(n235) );
  AOI33D0 U729 ( .A1(n321), .A2(port_dest[20]), .A3(port_dest[21]), .B1(n322), 
        .B2(port_dest[12]), .B3(port_dest[13]), .ZN(n320) );
  AOI33D0 U730 ( .A1(n323), .A2(port_dest[4]), .A3(port_dest[5]), .B1(n324), 
        .B2(port_dest[16]), .B3(port_dest[17]), .ZN(n319) );
  AOI33D0 U731 ( .A1(n325), .A2(port_dest[24]), .A3(port_dest[25]), .B1(n326), 
        .B2(port_dest[28]), .B3(port_dest[29]), .ZN(n318) );
  AOI33D0 U732 ( .A1(port_dest[0]), .A2(n327), .A3(n280), .B1(port_dest[8]), 
        .B2(n313), .B3(n103), .ZN(n317) );
  ND3D0 U733 ( .A1(n242), .A2(n244), .A3(n243), .ZN(n236) );
  ND3D0 U734 ( .A1(n37), .A2(n31), .A3(n34), .ZN(n316) );
  OAI21D0 U735 ( .A1(n43), .A2(port_dest[23]), .B(n328), .ZN(n34) );
  CKND2D0 U736 ( .A1(n43), .A2(port_dest[23]), .ZN(n37) );
  CKND0 U737 ( .I(n307), .ZN(n33) );
  CKND2D0 U738 ( .A1(n40), .A2(n212), .ZN(n307) );
  CKND2D0 U739 ( .A1(n41), .A2(n213), .ZN(n212) );
  NR2D0 U740 ( .A1(n328), .A2(n43), .ZN(n41) );
  AN2D0 U741 ( .A1(n29), .A2(port_dest[27]), .Z(n43) );
  OA21D0 U742 ( .A1(port_dest[27]), .A2(n29), .B(n329), .Z(n328) );
  NR2D0 U743 ( .A1(n81), .A2(n78), .ZN(n40) );
  NR2D0 U744 ( .A1(n21), .A2(port_dest[27]), .ZN(n78) );
  CKND0 U745 ( .I(n315), .ZN(n21) );
  NR2D0 U746 ( .A1(n329), .A2(n29), .ZN(n315) );
  NR2D0 U747 ( .A1(n244), .A2(n7), .ZN(n29) );
  AOI21D0 U748 ( .A1(n7), .A2(n244), .B(n242), .ZN(n329) );
  IND2D0 U749 ( .A1(n243), .B1(n234), .ZN(n81) );
  ND3D0 U750 ( .A1(n244), .A2(n7), .A3(n242), .ZN(n234) );
  ND4D0 U751 ( .A1(n330), .A2(n331), .A3(n332), .A4(n333), .ZN(n242) );
  AOI33D0 U752 ( .A1(port_dest[20]), .A2(n214), .A3(n321), .B1(port_dest[12]), 
        .B2(n304), .B3(n322), .ZN(n333) );
  AOI33D0 U753 ( .A1(port_dest[4]), .A2(n137), .A3(n323), .B1(port_dest[16]), 
        .B2(n303), .B3(n324), .ZN(n332) );
  AOI33D0 U754 ( .A1(port_dest[24]), .A2(n302), .A3(n325), .B1(port_dest[28]), 
        .B2(n229), .B3(n326), .ZN(n331) );
  AOI32D0 U755 ( .A1(n305), .A2(n327), .A3(port_dest[0]), .B1(n334), .B2(
        port_dest[8]), .ZN(n330) );
  ND4D0 U756 ( .A1(n335), .A2(n336), .A3(n337), .A4(n338), .ZN(n244) );
  AOI33D0 U757 ( .A1(n292), .A2(n214), .A3(n321), .B1(n294), .B2(n304), .B3(
        n322), .ZN(n338) );
  CKND0 U758 ( .I(port_dest[13]), .ZN(n304) );
  CKND0 U759 ( .I(port_dest[21]), .ZN(n214) );
  AOI33D0 U760 ( .A1(n290), .A2(n137), .A3(n323), .B1(n293), .B2(n303), .B3(
        n324), .ZN(n337) );
  CKND0 U761 ( .I(port_dest[17]), .ZN(n303) );
  CKND0 U762 ( .I(port_dest[5]), .ZN(n137) );
  AOI33D0 U763 ( .A1(n291), .A2(n302), .A3(n325), .B1(n289), .B2(n229), .B3(
        n326), .ZN(n336) );
  CKND0 U764 ( .I(port_dest[29]), .ZN(n229) );
  CKND0 U765 ( .I(port_dest[25]), .ZN(n302) );
  AOI32D0 U766 ( .A1(n146), .A2(n327), .A3(n305), .B1(n334), .B2(n295), .ZN(
        n335) );
  NR3D0 U767 ( .A1(port_dest[10]), .A2(port_dest[9]), .A3(n177), .ZN(n334) );
  NR2D0 U768 ( .A1(n100), .A2(port_dest[1]), .ZN(n305) );
  CKND0 U769 ( .I(port_dest[3]), .ZN(n100) );
  ND4D0 U770 ( .A1(n339), .A2(n340), .A3(n341), .A4(n342), .ZN(n243) );
  AOI33D0 U771 ( .A1(n321), .A2(n292), .A3(port_dest[21]), .B1(n322), .B2(n294), .B3(port_dest[13]), .ZN(n342) );
  CKND0 U772 ( .I(port_dest[12]), .ZN(n294) );
  NR2D0 U773 ( .A1(n248), .A2(port_dest[14]), .ZN(n322) );
  CKND0 U774 ( .I(port_dest[15]), .ZN(n248) );
  CKND0 U775 ( .I(port_dest[20]), .ZN(n292) );
  NR2D0 U776 ( .A1(n213), .A2(port_dest[22]), .ZN(n321) );
  CKND0 U777 ( .I(port_dest[23]), .ZN(n213) );
  AOI33D0 U778 ( .A1(n323), .A2(n290), .A3(port_dest[5]), .B1(n324), .B2(n293), 
        .B3(port_dest[17]), .ZN(n341) );
  CKND0 U779 ( .I(port_dest[16]), .ZN(n293) );
  NR2D0 U780 ( .A1(n31), .A2(port_dest[18]), .ZN(n324) );
  CKND0 U781 ( .I(port_dest[19]), .ZN(n31) );
  CKND0 U782 ( .I(port_dest[4]), .ZN(n290) );
  NR2D0 U783 ( .A1(n125), .A2(port_dest[6]), .ZN(n323) );
  CKND0 U784 ( .I(port_dest[7]), .ZN(n125) );
  AOI33D0 U785 ( .A1(n325), .A2(n291), .A3(port_dest[25]), .B1(n326), .B2(n289), .B3(port_dest[29]), .ZN(n340) );
  CKND0 U786 ( .I(port_dest[28]), .ZN(n289) );
  NR2D0 U787 ( .A1(n7), .A2(port_dest[30]), .ZN(n326) );
  CKND0 U788 ( .I(port_dest[31]), .ZN(n7) );
  CKND0 U789 ( .I(port_dest[24]), .ZN(n291) );
  NR2D0 U790 ( .A1(n19), .A2(port_dest[26]), .ZN(n325) );
  CKND0 U791 ( .I(port_dest[27]), .ZN(n19) );
  AOI33D0 U792 ( .A1(n146), .A2(n327), .A3(n280), .B1(n313), .B2(n295), .B3(
        n103), .ZN(n339) );
  NR2D0 U793 ( .A1(n301), .A2(n177), .ZN(n103) );
  CKND0 U794 ( .I(port_dest[11]), .ZN(n177) );
  CKND0 U795 ( .I(port_dest[9]), .ZN(n301) );
  CKND0 U796 ( .I(port_dest[8]), .ZN(n295) );
  CKND0 U797 ( .I(port_dest[10]), .ZN(n313) );
  CKND0 U798 ( .I(n96), .ZN(n280) );
  CKND2D0 U799 ( .A1(port_dest[1]), .A2(port_dest[3]), .ZN(n96) );
  CKND0 U800 ( .I(port_dest[2]), .ZN(n327) );
  CKND0 U801 ( .I(port_dest[0]), .ZN(n146) );
endmodule


module crossbar_0 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_1 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_2 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_3 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_4 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_5 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_6 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_7 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_8 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_9 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_10 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_11 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_12 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_13 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_14 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_15 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_16 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_17 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_18 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_19 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U82 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U83 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U84 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U85 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U86 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U87 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U88 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U89 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U90 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U91 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U92 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U93 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U94 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U95 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U96 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U97 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U98 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U99 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U100 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U101 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U102 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U103 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U104 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U105 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U106 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U107 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U108 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U109 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U110 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U111 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U112 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U113 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U114 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U115 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U116 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U117 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U118 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U119 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U120 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U121 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U122 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U123 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U124 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U125 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U126 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U127 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U128 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U129 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U130 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U131 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U132 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U133 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U134 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U135 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U136 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U137 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U138 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U139 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U140 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U141 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U142 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U143 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U144 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U145 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U146 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U147 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U148 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U149 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U150 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U151 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U152 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U153 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U154 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U155 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U156 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U157 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U158 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U159 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U160 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U161 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module benes ( in_input, in_control, port_en_n, out_output, clk, rst );
  input [127:0] in_input;
  input [19:0] in_control;
  input [7:0] port_en_n;
  output [159:0] out_output;
  input clk, rst;
  wire   \*Logic1* , \in_upper_00[3] , \in_lower_00[3] , \in_upper_01[3] ,
         \in_lower_01[3] , in_upper_02_3, \in_lower_02[3] , \in_upper_03[3] ,
         \stage_0_output[7][19] , \stage_0_output[7][18] ,
         \stage_0_output[7][17] , \stage_0_output[7][16] ,
         \stage_0_output[7][15] , \stage_0_output[7][14] ,
         \stage_0_output[7][13] , \stage_0_output[7][12] ,
         \stage_0_output[7][11] , \stage_0_output[7][10] ,
         \stage_0_output[7][9] , \stage_0_output[7][8] ,
         \stage_0_output[7][7] , \stage_0_output[7][6] ,
         \stage_0_output[7][5] , \stage_0_output[7][4] ,
         \stage_0_output[7][3] , \stage_0_output[7][2] ,
         \stage_0_output[7][1] , \stage_0_output[7][0] ,
         \stage_0_output[6][19] , \stage_0_output[6][18] ,
         \stage_0_output[6][17] , \stage_0_output[6][16] ,
         \stage_0_output[6][15] , \stage_0_output[6][14] ,
         \stage_0_output[6][13] , \stage_0_output[6][12] ,
         \stage_0_output[6][11] , \stage_0_output[6][10] ,
         \stage_0_output[6][9] , \stage_0_output[6][8] ,
         \stage_0_output[6][7] , \stage_0_output[6][6] ,
         \stage_0_output[6][5] , \stage_0_output[6][4] ,
         \stage_0_output[6][3] , \stage_0_output[6][2] ,
         \stage_0_output[6][1] , \stage_0_output[6][0] ,
         \stage_0_output[5][19] , \stage_0_output[5][18] ,
         \stage_0_output[5][17] , \stage_0_output[5][16] ,
         \stage_0_output[5][15] , \stage_0_output[5][14] ,
         \stage_0_output[5][13] , \stage_0_output[5][12] ,
         \stage_0_output[5][11] , \stage_0_output[5][10] ,
         \stage_0_output[5][9] , \stage_0_output[5][8] ,
         \stage_0_output[5][7] , \stage_0_output[5][6] ,
         \stage_0_output[5][5] , \stage_0_output[5][4] ,
         \stage_0_output[5][3] , \stage_0_output[5][2] ,
         \stage_0_output[5][1] , \stage_0_output[5][0] ,
         \stage_0_output[4][19] , \stage_0_output[4][18] ,
         \stage_0_output[4][17] , \stage_0_output[4][16] ,
         \stage_0_output[4][15] , \stage_0_output[4][14] ,
         \stage_0_output[4][13] , \stage_0_output[4][12] ,
         \stage_0_output[4][11] , \stage_0_output[4][10] ,
         \stage_0_output[4][9] , \stage_0_output[4][8] ,
         \stage_0_output[4][7] , \stage_0_output[4][6] ,
         \stage_0_output[4][5] , \stage_0_output[4][4] ,
         \stage_0_output[4][3] , \stage_0_output[4][2] ,
         \stage_0_output[4][1] , \stage_0_output[4][0] ,
         \stage_0_output[3][19] , \stage_0_output[3][18] ,
         \stage_0_output[3][17] , \stage_0_output[3][16] ,
         \stage_0_output[3][15] , \stage_0_output[3][14] ,
         \stage_0_output[3][13] , \stage_0_output[3][12] ,
         \stage_0_output[3][11] , \stage_0_output[3][10] ,
         \stage_0_output[3][9] , \stage_0_output[3][8] ,
         \stage_0_output[3][7] , \stage_0_output[3][6] ,
         \stage_0_output[3][5] , \stage_0_output[3][4] ,
         \stage_0_output[3][3] , \stage_0_output[3][2] ,
         \stage_0_output[3][1] , \stage_0_output[3][0] ,
         \stage_0_output[2][19] , \stage_0_output[2][18] ,
         \stage_0_output[2][17] , \stage_0_output[2][16] ,
         \stage_0_output[2][15] , \stage_0_output[2][14] ,
         \stage_0_output[2][13] , \stage_0_output[2][12] ,
         \stage_0_output[2][11] , \stage_0_output[2][10] ,
         \stage_0_output[2][9] , \stage_0_output[2][8] ,
         \stage_0_output[2][7] , \stage_0_output[2][6] ,
         \stage_0_output[2][5] , \stage_0_output[2][4] ,
         \stage_0_output[2][3] , \stage_0_output[2][2] ,
         \stage_0_output[2][1] , \stage_0_output[2][0] ,
         \stage_0_output[1][19] , \stage_0_output[1][18] ,
         \stage_0_output[1][17] , \stage_0_output[1][16] ,
         \stage_0_output[1][15] , \stage_0_output[1][14] ,
         \stage_0_output[1][13] , \stage_0_output[1][12] ,
         \stage_0_output[1][11] , \stage_0_output[1][10] ,
         \stage_0_output[1][9] , \stage_0_output[1][8] ,
         \stage_0_output[1][7] , \stage_0_output[1][6] ,
         \stage_0_output[1][5] , \stage_0_output[1][4] ,
         \stage_0_output[1][3] , \stage_0_output[1][2] ,
         \stage_0_output[1][1] , \stage_0_output[1][0] ,
         \stage_0_output[0][19] , \stage_0_output[0][18] ,
         \stage_0_output[0][17] , \stage_0_output[0][16] ,
         \stage_0_output[0][15] , \stage_0_output[0][14] ,
         \stage_0_output[0][13] , \stage_0_output[0][12] ,
         \stage_0_output[0][11] , \stage_0_output[0][10] ,
         \stage_0_output[0][9] , \stage_0_output[0][8] ,
         \stage_0_output[0][7] , \stage_0_output[0][6] ,
         \stage_0_output[0][5] , \stage_0_output[0][4] ,
         \stage_0_output[0][3] , \stage_0_output[0][2] ,
         \stage_0_output[0][1] , \stage_0_output[0][0] ,
         \stage_0_retimer[7][19] , \stage_0_retimer[7][18] ,
         \stage_0_retimer[7][17] , \stage_0_retimer[7][16] ,
         \stage_0_retimer[7][15] , \stage_0_retimer[7][14] ,
         \stage_0_retimer[7][13] , \stage_0_retimer[7][12] ,
         \stage_0_retimer[7][11] , \stage_0_retimer[7][10] ,
         \stage_0_retimer[7][9] , \stage_0_retimer[7][8] ,
         \stage_0_retimer[7][7] , \stage_0_retimer[7][6] ,
         \stage_0_retimer[7][5] , \stage_0_retimer[7][4] ,
         \stage_0_retimer[7][3] , \stage_0_retimer[7][2] ,
         \stage_0_retimer[7][1] , \stage_0_retimer[7][0] ,
         \stage_0_retimer[6][19] , \stage_0_retimer[6][18] ,
         \stage_0_retimer[6][17] , \stage_0_retimer[6][16] ,
         \stage_0_retimer[6][15] , \stage_0_retimer[6][14] ,
         \stage_0_retimer[6][13] , \stage_0_retimer[6][12] ,
         \stage_0_retimer[6][11] , \stage_0_retimer[6][10] ,
         \stage_0_retimer[6][9] , \stage_0_retimer[6][8] ,
         \stage_0_retimer[6][7] , \stage_0_retimer[6][6] ,
         \stage_0_retimer[6][5] , \stage_0_retimer[6][4] ,
         \stage_0_retimer[6][3] , \stage_0_retimer[6][2] ,
         \stage_0_retimer[6][1] , \stage_0_retimer[6][0] ,
         \stage_0_retimer[5][19] , \stage_0_retimer[5][18] ,
         \stage_0_retimer[5][17] , \stage_0_retimer[5][16] ,
         \stage_0_retimer[5][15] , \stage_0_retimer[5][14] ,
         \stage_0_retimer[5][13] , \stage_0_retimer[5][12] ,
         \stage_0_retimer[5][11] , \stage_0_retimer[5][10] ,
         \stage_0_retimer[5][9] , \stage_0_retimer[5][8] ,
         \stage_0_retimer[5][7] , \stage_0_retimer[5][6] ,
         \stage_0_retimer[5][5] , \stage_0_retimer[5][4] ,
         \stage_0_retimer[5][3] , \stage_0_retimer[5][2] ,
         \stage_0_retimer[5][1] , \stage_0_retimer[5][0] ,
         \stage_0_retimer[4][19] , \stage_0_retimer[4][18] ,
         \stage_0_retimer[4][17] , \stage_0_retimer[4][16] ,
         \stage_0_retimer[4][15] , \stage_0_retimer[4][14] ,
         \stage_0_retimer[4][13] , \stage_0_retimer[4][12] ,
         \stage_0_retimer[4][11] , \stage_0_retimer[4][10] ,
         \stage_0_retimer[4][9] , \stage_0_retimer[4][8] ,
         \stage_0_retimer[4][7] , \stage_0_retimer[4][6] ,
         \stage_0_retimer[4][5] , \stage_0_retimer[4][4] ,
         \stage_0_retimer[4][3] , \stage_0_retimer[4][2] ,
         \stage_0_retimer[4][1] , \stage_0_retimer[4][0] ,
         \stage_0_retimer[3][19] , \stage_0_retimer[3][18] ,
         \stage_0_retimer[3][17] , \stage_0_retimer[3][16] ,
         \stage_0_retimer[3][15] , \stage_0_retimer[3][14] ,
         \stage_0_retimer[3][13] , \stage_0_retimer[3][12] ,
         \stage_0_retimer[3][11] , \stage_0_retimer[3][10] ,
         \stage_0_retimer[3][9] , \stage_0_retimer[3][8] ,
         \stage_0_retimer[3][7] , \stage_0_retimer[3][6] ,
         \stage_0_retimer[3][5] , \stage_0_retimer[3][4] ,
         \stage_0_retimer[3][3] , \stage_0_retimer[3][2] ,
         \stage_0_retimer[3][1] , \stage_0_retimer[3][0] ,
         \stage_0_retimer[2][19] , \stage_0_retimer[2][18] ,
         \stage_0_retimer[2][17] , \stage_0_retimer[2][16] ,
         \stage_0_retimer[2][15] , \stage_0_retimer[2][14] ,
         \stage_0_retimer[2][13] , \stage_0_retimer[2][12] ,
         \stage_0_retimer[2][11] , \stage_0_retimer[2][10] ,
         \stage_0_retimer[2][9] , \stage_0_retimer[2][8] ,
         \stage_0_retimer[2][7] , \stage_0_retimer[2][6] ,
         \stage_0_retimer[2][5] , \stage_0_retimer[2][4] ,
         \stage_0_retimer[2][3] , \stage_0_retimer[2][2] ,
         \stage_0_retimer[2][1] , \stage_0_retimer[2][0] ,
         \stage_0_retimer[1][19] , \stage_0_retimer[1][18] ,
         \stage_0_retimer[1][17] , \stage_0_retimer[1][16] ,
         \stage_0_retimer[1][15] , \stage_0_retimer[1][14] ,
         \stage_0_retimer[1][13] , \stage_0_retimer[1][12] ,
         \stage_0_retimer[1][11] , \stage_0_retimer[1][10] ,
         \stage_0_retimer[1][9] , \stage_0_retimer[1][8] ,
         \stage_0_retimer[1][7] , \stage_0_retimer[1][6] ,
         \stage_0_retimer[1][5] , \stage_0_retimer[1][4] ,
         \stage_0_retimer[1][3] , \stage_0_retimer[1][2] ,
         \stage_0_retimer[1][1] , \stage_0_retimer[1][0] ,
         \stage_0_retimer[0][19] , \stage_0_retimer[0][18] ,
         \stage_0_retimer[0][17] , \stage_0_retimer[0][16] ,
         \stage_0_retimer[0][15] , \stage_0_retimer[0][14] ,
         \stage_0_retimer[0][13] , \stage_0_retimer[0][12] ,
         \stage_0_retimer[0][11] , \stage_0_retimer[0][10] ,
         \stage_0_retimer[0][9] , \stage_0_retimer[0][8] ,
         \stage_0_retimer[0][7] , \stage_0_retimer[0][6] ,
         \stage_0_retimer[0][5] , \stage_0_retimer[0][4] ,
         \stage_0_retimer[0][3] , \stage_0_retimer[0][2] ,
         \stage_0_retimer[0][1] , \stage_0_retimer[0][0] ,
         \stage_1_output[7][19] , \stage_1_output[7][18] ,
         \stage_1_output[7][17] , \stage_1_output[7][16] ,
         \stage_1_output[7][15] , \stage_1_output[7][14] ,
         \stage_1_output[7][13] , \stage_1_output[7][12] ,
         \stage_1_output[7][11] , \stage_1_output[7][10] ,
         \stage_1_output[7][9] , \stage_1_output[7][8] ,
         \stage_1_output[7][7] , \stage_1_output[7][6] ,
         \stage_1_output[7][5] , \stage_1_output[7][4] ,
         \stage_1_output[7][3] , \stage_1_output[7][2] ,
         \stage_1_output[7][1] , \stage_1_output[7][0] ,
         \stage_1_output[6][19] , \stage_1_output[6][18] ,
         \stage_1_output[6][17] , \stage_1_output[6][16] ,
         \stage_1_output[6][15] , \stage_1_output[6][14] ,
         \stage_1_output[6][13] , \stage_1_output[6][12] ,
         \stage_1_output[6][11] , \stage_1_output[6][10] ,
         \stage_1_output[6][9] , \stage_1_output[6][8] ,
         \stage_1_output[6][7] , \stage_1_output[6][6] ,
         \stage_1_output[6][5] , \stage_1_output[6][4] ,
         \stage_1_output[6][3] , \stage_1_output[6][2] ,
         \stage_1_output[6][1] , \stage_1_output[6][0] ,
         \stage_1_output[5][19] , \stage_1_output[5][18] ,
         \stage_1_output[5][17] , \stage_1_output[5][16] ,
         \stage_1_output[5][15] , \stage_1_output[5][14] ,
         \stage_1_output[5][13] , \stage_1_output[5][12] ,
         \stage_1_output[5][11] , \stage_1_output[5][10] ,
         \stage_1_output[5][9] , \stage_1_output[5][8] ,
         \stage_1_output[5][7] , \stage_1_output[5][6] ,
         \stage_1_output[5][5] , \stage_1_output[5][4] ,
         \stage_1_output[5][3] , \stage_1_output[5][2] ,
         \stage_1_output[5][1] , \stage_1_output[5][0] ,
         \stage_1_output[4][19] , \stage_1_output[4][18] ,
         \stage_1_output[4][17] , \stage_1_output[4][16] ,
         \stage_1_output[4][15] , \stage_1_output[4][14] ,
         \stage_1_output[4][13] , \stage_1_output[4][12] ,
         \stage_1_output[4][11] , \stage_1_output[4][10] ,
         \stage_1_output[4][9] , \stage_1_output[4][8] ,
         \stage_1_output[4][7] , \stage_1_output[4][6] ,
         \stage_1_output[4][5] , \stage_1_output[4][4] ,
         \stage_1_output[4][3] , \stage_1_output[4][2] ,
         \stage_1_output[4][1] , \stage_1_output[4][0] ,
         \stage_1_output[3][19] , \stage_1_output[3][18] ,
         \stage_1_output[3][17] , \stage_1_output[3][16] ,
         \stage_1_output[3][15] , \stage_1_output[3][14] ,
         \stage_1_output[3][13] , \stage_1_output[3][12] ,
         \stage_1_output[3][11] , \stage_1_output[3][10] ,
         \stage_1_output[3][9] , \stage_1_output[3][8] ,
         \stage_1_output[3][7] , \stage_1_output[3][6] ,
         \stage_1_output[3][5] , \stage_1_output[3][4] ,
         \stage_1_output[3][3] , \stage_1_output[3][2] ,
         \stage_1_output[3][1] , \stage_1_output[3][0] ,
         \stage_1_output[2][19] , \stage_1_output[2][18] ,
         \stage_1_output[2][17] , \stage_1_output[2][16] ,
         \stage_1_output[2][15] , \stage_1_output[2][14] ,
         \stage_1_output[2][13] , \stage_1_output[2][12] ,
         \stage_1_output[2][11] , \stage_1_output[2][10] ,
         \stage_1_output[2][9] , \stage_1_output[2][8] ,
         \stage_1_output[2][7] , \stage_1_output[2][6] ,
         \stage_1_output[2][5] , \stage_1_output[2][4] ,
         \stage_1_output[2][3] , \stage_1_output[2][2] ,
         \stage_1_output[2][1] , \stage_1_output[2][0] ,
         \stage_1_output[1][19] , \stage_1_output[1][18] ,
         \stage_1_output[1][17] , \stage_1_output[1][16] ,
         \stage_1_output[1][15] , \stage_1_output[1][14] ,
         \stage_1_output[1][13] , \stage_1_output[1][12] ,
         \stage_1_output[1][11] , \stage_1_output[1][10] ,
         \stage_1_output[1][9] , \stage_1_output[1][8] ,
         \stage_1_output[1][7] , \stage_1_output[1][6] ,
         \stage_1_output[1][5] , \stage_1_output[1][4] ,
         \stage_1_output[1][3] , \stage_1_output[1][2] ,
         \stage_1_output[1][1] , \stage_1_output[1][0] ,
         \stage_1_output[0][19] , \stage_1_output[0][18] ,
         \stage_1_output[0][17] , \stage_1_output[0][16] ,
         \stage_1_output[0][15] , \stage_1_output[0][14] ,
         \stage_1_output[0][13] , \stage_1_output[0][12] ,
         \stage_1_output[0][11] , \stage_1_output[0][10] ,
         \stage_1_output[0][9] , \stage_1_output[0][8] ,
         \stage_1_output[0][7] , \stage_1_output[0][6] ,
         \stage_1_output[0][5] , \stage_1_output[0][4] ,
         \stage_1_output[0][3] , \stage_1_output[0][2] ,
         \stage_1_output[0][1] , \stage_1_output[0][0] ,
         \stage_1_retimer[7][19] , \stage_1_retimer[7][18] ,
         \stage_1_retimer[7][17] , \stage_1_retimer[7][16] ,
         \stage_1_retimer[7][15] , \stage_1_retimer[7][14] ,
         \stage_1_retimer[7][13] , \stage_1_retimer[7][12] ,
         \stage_1_retimer[7][11] , \stage_1_retimer[7][10] ,
         \stage_1_retimer[7][9] , \stage_1_retimer[7][8] ,
         \stage_1_retimer[7][7] , \stage_1_retimer[7][6] ,
         \stage_1_retimer[7][5] , \stage_1_retimer[7][4] ,
         \stage_1_retimer[7][3] , \stage_1_retimer[7][2] ,
         \stage_1_retimer[7][1] , \stage_1_retimer[7][0] ,
         \stage_1_retimer[6][19] , \stage_1_retimer[6][18] ,
         \stage_1_retimer[6][17] , \stage_1_retimer[6][16] ,
         \stage_1_retimer[6][15] , \stage_1_retimer[6][14] ,
         \stage_1_retimer[6][13] , \stage_1_retimer[6][12] ,
         \stage_1_retimer[6][11] , \stage_1_retimer[6][10] ,
         \stage_1_retimer[6][9] , \stage_1_retimer[6][8] ,
         \stage_1_retimer[6][7] , \stage_1_retimer[6][6] ,
         \stage_1_retimer[6][5] , \stage_1_retimer[6][4] ,
         \stage_1_retimer[6][3] , \stage_1_retimer[6][2] ,
         \stage_1_retimer[6][1] , \stage_1_retimer[6][0] ,
         \stage_1_retimer[5][19] , \stage_1_retimer[5][18] ,
         \stage_1_retimer[5][17] , \stage_1_retimer[5][16] ,
         \stage_1_retimer[5][15] , \stage_1_retimer[5][14] ,
         \stage_1_retimer[5][13] , \stage_1_retimer[5][12] ,
         \stage_1_retimer[5][11] , \stage_1_retimer[5][10] ,
         \stage_1_retimer[5][9] , \stage_1_retimer[5][8] ,
         \stage_1_retimer[5][7] , \stage_1_retimer[5][6] ,
         \stage_1_retimer[5][5] , \stage_1_retimer[5][4] ,
         \stage_1_retimer[5][3] , \stage_1_retimer[5][2] ,
         \stage_1_retimer[5][1] , \stage_1_retimer[5][0] ,
         \stage_1_retimer[4][19] , \stage_1_retimer[4][18] ,
         \stage_1_retimer[4][17] , \stage_1_retimer[4][16] ,
         \stage_1_retimer[4][15] , \stage_1_retimer[4][14] ,
         \stage_1_retimer[4][13] , \stage_1_retimer[4][12] ,
         \stage_1_retimer[4][11] , \stage_1_retimer[4][10] ,
         \stage_1_retimer[4][9] , \stage_1_retimer[4][8] ,
         \stage_1_retimer[4][7] , \stage_1_retimer[4][6] ,
         \stage_1_retimer[4][5] , \stage_1_retimer[4][4] ,
         \stage_1_retimer[4][3] , \stage_1_retimer[4][2] ,
         \stage_1_retimer[4][1] , \stage_1_retimer[4][0] ,
         \stage_1_retimer[3][19] , \stage_1_retimer[3][18] ,
         \stage_1_retimer[3][17] , \stage_1_retimer[3][16] ,
         \stage_1_retimer[3][15] , \stage_1_retimer[3][14] ,
         \stage_1_retimer[3][13] , \stage_1_retimer[3][12] ,
         \stage_1_retimer[3][11] , \stage_1_retimer[3][10] ,
         \stage_1_retimer[3][9] , \stage_1_retimer[3][8] ,
         \stage_1_retimer[3][7] , \stage_1_retimer[3][6] ,
         \stage_1_retimer[3][5] , \stage_1_retimer[3][4] ,
         \stage_1_retimer[3][3] , \stage_1_retimer[3][2] ,
         \stage_1_retimer[3][1] , \stage_1_retimer[3][0] ,
         \stage_1_retimer[2][19] , \stage_1_retimer[2][18] ,
         \stage_1_retimer[2][17] , \stage_1_retimer[2][16] ,
         \stage_1_retimer[2][15] , \stage_1_retimer[2][14] ,
         \stage_1_retimer[2][13] , \stage_1_retimer[2][12] ,
         \stage_1_retimer[2][11] , \stage_1_retimer[2][10] ,
         \stage_1_retimer[2][9] , \stage_1_retimer[2][8] ,
         \stage_1_retimer[2][7] , \stage_1_retimer[2][6] ,
         \stage_1_retimer[2][5] , \stage_1_retimer[2][4] ,
         \stage_1_retimer[2][3] , \stage_1_retimer[2][2] ,
         \stage_1_retimer[2][1] , \stage_1_retimer[2][0] ,
         \stage_1_retimer[1][19] , \stage_1_retimer[1][18] ,
         \stage_1_retimer[1][17] , \stage_1_retimer[1][16] ,
         \stage_1_retimer[1][15] , \stage_1_retimer[1][14] ,
         \stage_1_retimer[1][13] , \stage_1_retimer[1][12] ,
         \stage_1_retimer[1][11] , \stage_1_retimer[1][10] ,
         \stage_1_retimer[1][9] , \stage_1_retimer[1][8] ,
         \stage_1_retimer[1][7] , \stage_1_retimer[1][6] ,
         \stage_1_retimer[1][5] , \stage_1_retimer[1][4] ,
         \stage_1_retimer[1][3] , \stage_1_retimer[1][2] ,
         \stage_1_retimer[1][1] , \stage_1_retimer[1][0] ,
         \stage_1_retimer[0][19] , \stage_1_retimer[0][18] ,
         \stage_1_retimer[0][17] , \stage_1_retimer[0][16] ,
         \stage_1_retimer[0][15] , \stage_1_retimer[0][14] ,
         \stage_1_retimer[0][13] , \stage_1_retimer[0][12] ,
         \stage_1_retimer[0][11] , \stage_1_retimer[0][10] ,
         \stage_1_retimer[0][9] , \stage_1_retimer[0][8] ,
         \stage_1_retimer[0][7] , \stage_1_retimer[0][6] ,
         \stage_1_retimer[0][5] , \stage_1_retimer[0][4] ,
         \stage_1_retimer[0][3] , \stage_1_retimer[0][2] ,
         \stage_1_retimer[0][1] , \stage_1_retimer[0][0] ,
         \stage_2_output[7][19] , \stage_2_output[7][18] ,
         \stage_2_output[7][17] , \stage_2_output[7][16] ,
         \stage_2_output[7][15] , \stage_2_output[7][14] ,
         \stage_2_output[7][13] , \stage_2_output[7][12] ,
         \stage_2_output[7][11] , \stage_2_output[7][10] ,
         \stage_2_output[7][9] , \stage_2_output[7][8] ,
         \stage_2_output[7][7] , \stage_2_output[7][6] ,
         \stage_2_output[7][5] , \stage_2_output[7][4] ,
         \stage_2_output[7][3] , \stage_2_output[7][2] ,
         \stage_2_output[7][1] , \stage_2_output[7][0] ,
         \stage_2_output[6][19] , \stage_2_output[6][18] ,
         \stage_2_output[6][17] , \stage_2_output[6][16] ,
         \stage_2_output[6][15] , \stage_2_output[6][14] ,
         \stage_2_output[6][13] , \stage_2_output[6][12] ,
         \stage_2_output[6][11] , \stage_2_output[6][10] ,
         \stage_2_output[6][9] , \stage_2_output[6][8] ,
         \stage_2_output[6][7] , \stage_2_output[6][6] ,
         \stage_2_output[6][5] , \stage_2_output[6][4] ,
         \stage_2_output[6][3] , \stage_2_output[6][2] ,
         \stage_2_output[6][1] , \stage_2_output[6][0] ,
         \stage_2_output[5][19] , \stage_2_output[5][18] ,
         \stage_2_output[5][17] , \stage_2_output[5][16] ,
         \stage_2_output[5][15] , \stage_2_output[5][14] ,
         \stage_2_output[5][13] , \stage_2_output[5][12] ,
         \stage_2_output[5][11] , \stage_2_output[5][10] ,
         \stage_2_output[5][9] , \stage_2_output[5][8] ,
         \stage_2_output[5][7] , \stage_2_output[5][6] ,
         \stage_2_output[5][5] , \stage_2_output[5][4] ,
         \stage_2_output[5][3] , \stage_2_output[5][2] ,
         \stage_2_output[5][1] , \stage_2_output[5][0] ,
         \stage_2_output[4][19] , \stage_2_output[4][18] ,
         \stage_2_output[4][17] , \stage_2_output[4][16] ,
         \stage_2_output[4][15] , \stage_2_output[4][14] ,
         \stage_2_output[4][13] , \stage_2_output[4][12] ,
         \stage_2_output[4][11] , \stage_2_output[4][10] ,
         \stage_2_output[4][9] , \stage_2_output[4][8] ,
         \stage_2_output[4][7] , \stage_2_output[4][6] ,
         \stage_2_output[4][5] , \stage_2_output[4][4] ,
         \stage_2_output[4][3] , \stage_2_output[4][2] ,
         \stage_2_output[4][1] , \stage_2_output[4][0] ,
         \stage_2_output[3][19] , \stage_2_output[3][18] ,
         \stage_2_output[3][17] , \stage_2_output[3][16] ,
         \stage_2_output[3][15] , \stage_2_output[3][14] ,
         \stage_2_output[3][13] , \stage_2_output[3][12] ,
         \stage_2_output[3][11] , \stage_2_output[3][10] ,
         \stage_2_output[3][9] , \stage_2_output[3][8] ,
         \stage_2_output[3][7] , \stage_2_output[3][6] ,
         \stage_2_output[3][5] , \stage_2_output[3][4] ,
         \stage_2_output[3][3] , \stage_2_output[3][2] ,
         \stage_2_output[3][1] , \stage_2_output[3][0] ,
         \stage_2_output[2][19] , \stage_2_output[2][18] ,
         \stage_2_output[2][17] , \stage_2_output[2][16] ,
         \stage_2_output[2][15] , \stage_2_output[2][14] ,
         \stage_2_output[2][13] , \stage_2_output[2][12] ,
         \stage_2_output[2][11] , \stage_2_output[2][10] ,
         \stage_2_output[2][9] , \stage_2_output[2][8] ,
         \stage_2_output[2][7] , \stage_2_output[2][6] ,
         \stage_2_output[2][5] , \stage_2_output[2][4] ,
         \stage_2_output[2][3] , \stage_2_output[2][2] ,
         \stage_2_output[2][1] , \stage_2_output[2][0] ,
         \stage_2_output[1][19] , \stage_2_output[1][18] ,
         \stage_2_output[1][17] , \stage_2_output[1][16] ,
         \stage_2_output[1][15] , \stage_2_output[1][14] ,
         \stage_2_output[1][13] , \stage_2_output[1][12] ,
         \stage_2_output[1][11] , \stage_2_output[1][10] ,
         \stage_2_output[1][9] , \stage_2_output[1][8] ,
         \stage_2_output[1][7] , \stage_2_output[1][6] ,
         \stage_2_output[1][5] , \stage_2_output[1][4] ,
         \stage_2_output[1][3] , \stage_2_output[1][2] ,
         \stage_2_output[1][1] , \stage_2_output[1][0] ,
         \stage_2_output[0][19] , \stage_2_output[0][18] ,
         \stage_2_output[0][17] , \stage_2_output[0][16] ,
         \stage_2_output[0][15] , \stage_2_output[0][14] ,
         \stage_2_output[0][13] , \stage_2_output[0][12] ,
         \stage_2_output[0][11] , \stage_2_output[0][10] ,
         \stage_2_output[0][9] , \stage_2_output[0][8] ,
         \stage_2_output[0][7] , \stage_2_output[0][6] ,
         \stage_2_output[0][5] , \stage_2_output[0][4] ,
         \stage_2_output[0][3] , \stage_2_output[0][2] ,
         \stage_2_output[0][1] , \stage_2_output[0][0] ,
         \stage_2_retimer[7][19] , \stage_2_retimer[7][18] ,
         \stage_2_retimer[7][17] , \stage_2_retimer[7][16] ,
         \stage_2_retimer[7][15] , \stage_2_retimer[7][14] ,
         \stage_2_retimer[7][13] , \stage_2_retimer[7][12] ,
         \stage_2_retimer[7][11] , \stage_2_retimer[7][10] ,
         \stage_2_retimer[7][9] , \stage_2_retimer[7][8] ,
         \stage_2_retimer[7][7] , \stage_2_retimer[7][6] ,
         \stage_2_retimer[7][5] , \stage_2_retimer[7][4] ,
         \stage_2_retimer[7][3] , \stage_2_retimer[7][2] ,
         \stage_2_retimer[7][1] , \stage_2_retimer[7][0] ,
         \stage_2_retimer[6][19] , \stage_2_retimer[6][18] ,
         \stage_2_retimer[6][17] , \stage_2_retimer[6][16] ,
         \stage_2_retimer[6][15] , \stage_2_retimer[6][14] ,
         \stage_2_retimer[6][13] , \stage_2_retimer[6][12] ,
         \stage_2_retimer[6][11] , \stage_2_retimer[6][10] ,
         \stage_2_retimer[6][9] , \stage_2_retimer[6][8] ,
         \stage_2_retimer[6][7] , \stage_2_retimer[6][6] ,
         \stage_2_retimer[6][5] , \stage_2_retimer[6][4] ,
         \stage_2_retimer[6][3] , \stage_2_retimer[6][2] ,
         \stage_2_retimer[6][1] , \stage_2_retimer[6][0] ,
         \stage_2_retimer[5][19] , \stage_2_retimer[5][18] ,
         \stage_2_retimer[5][17] , \stage_2_retimer[5][16] ,
         \stage_2_retimer[5][15] , \stage_2_retimer[5][14] ,
         \stage_2_retimer[5][13] , \stage_2_retimer[5][12] ,
         \stage_2_retimer[5][11] , \stage_2_retimer[5][10] ,
         \stage_2_retimer[5][9] , \stage_2_retimer[5][8] ,
         \stage_2_retimer[5][7] , \stage_2_retimer[5][6] ,
         \stage_2_retimer[5][5] , \stage_2_retimer[5][4] ,
         \stage_2_retimer[5][3] , \stage_2_retimer[5][2] ,
         \stage_2_retimer[5][1] , \stage_2_retimer[5][0] ,
         \stage_2_retimer[4][19] , \stage_2_retimer[4][18] ,
         \stage_2_retimer[4][17] , \stage_2_retimer[4][16] ,
         \stage_2_retimer[4][15] , \stage_2_retimer[4][14] ,
         \stage_2_retimer[4][13] , \stage_2_retimer[4][12] ,
         \stage_2_retimer[4][11] , \stage_2_retimer[4][10] ,
         \stage_2_retimer[4][9] , \stage_2_retimer[4][8] ,
         \stage_2_retimer[4][7] , \stage_2_retimer[4][6] ,
         \stage_2_retimer[4][5] , \stage_2_retimer[4][4] ,
         \stage_2_retimer[4][3] , \stage_2_retimer[4][2] ,
         \stage_2_retimer[4][1] , \stage_2_retimer[4][0] ,
         \stage_2_retimer[3][19] , \stage_2_retimer[3][18] ,
         \stage_2_retimer[3][17] , \stage_2_retimer[3][16] ,
         \stage_2_retimer[3][15] , \stage_2_retimer[3][14] ,
         \stage_2_retimer[3][13] , \stage_2_retimer[3][12] ,
         \stage_2_retimer[3][11] , \stage_2_retimer[3][10] ,
         \stage_2_retimer[3][9] , \stage_2_retimer[3][8] ,
         \stage_2_retimer[3][7] , \stage_2_retimer[3][6] ,
         \stage_2_retimer[3][5] , \stage_2_retimer[3][4] ,
         \stage_2_retimer[3][3] , \stage_2_retimer[3][2] ,
         \stage_2_retimer[3][1] , \stage_2_retimer[3][0] ,
         \stage_2_retimer[2][19] , \stage_2_retimer[2][18] ,
         \stage_2_retimer[2][17] , \stage_2_retimer[2][16] ,
         \stage_2_retimer[2][15] , \stage_2_retimer[2][14] ,
         \stage_2_retimer[2][13] , \stage_2_retimer[2][12] ,
         \stage_2_retimer[2][11] , \stage_2_retimer[2][10] ,
         \stage_2_retimer[2][9] , \stage_2_retimer[2][8] ,
         \stage_2_retimer[2][7] , \stage_2_retimer[2][6] ,
         \stage_2_retimer[2][5] , \stage_2_retimer[2][4] ,
         \stage_2_retimer[2][3] , \stage_2_retimer[2][2] ,
         \stage_2_retimer[2][1] , \stage_2_retimer[2][0] ,
         \stage_2_retimer[1][19] , \stage_2_retimer[1][18] ,
         \stage_2_retimer[1][17] , \stage_2_retimer[1][16] ,
         \stage_2_retimer[1][15] , \stage_2_retimer[1][14] ,
         \stage_2_retimer[1][13] , \stage_2_retimer[1][12] ,
         \stage_2_retimer[1][11] , \stage_2_retimer[1][10] ,
         \stage_2_retimer[1][9] , \stage_2_retimer[1][8] ,
         \stage_2_retimer[1][7] , \stage_2_retimer[1][6] ,
         \stage_2_retimer[1][5] , \stage_2_retimer[1][4] ,
         \stage_2_retimer[1][3] , \stage_2_retimer[1][2] ,
         \stage_2_retimer[1][1] , \stage_2_retimer[1][0] ,
         \stage_2_retimer[0][19] , \stage_2_retimer[0][18] ,
         \stage_2_retimer[0][17] , \stage_2_retimer[0][16] ,
         \stage_2_retimer[0][15] , \stage_2_retimer[0][14] ,
         \stage_2_retimer[0][13] , \stage_2_retimer[0][12] ,
         \stage_2_retimer[0][11] , \stage_2_retimer[0][10] ,
         \stage_2_retimer[0][9] , \stage_2_retimer[0][8] ,
         \stage_2_retimer[0][7] , \stage_2_retimer[0][6] ,
         \stage_2_retimer[0][5] , \stage_2_retimer[0][4] ,
         \stage_2_retimer[0][3] , \stage_2_retimer[0][2] ,
         \stage_2_retimer[0][1] , \stage_2_retimer[0][0] ,
         \stage_3_output[7][19] , \stage_3_output[7][18] ,
         \stage_3_output[7][17] , \stage_3_output[7][16] ,
         \stage_3_output[7][15] , \stage_3_output[7][14] ,
         \stage_3_output[7][13] , \stage_3_output[7][12] ,
         \stage_3_output[7][11] , \stage_3_output[7][10] ,
         \stage_3_output[7][9] , \stage_3_output[7][8] ,
         \stage_3_output[7][7] , \stage_3_output[7][6] ,
         \stage_3_output[7][5] , \stage_3_output[7][4] ,
         \stage_3_output[7][3] , \stage_3_output[7][2] ,
         \stage_3_output[7][1] , \stage_3_output[7][0] ,
         \stage_3_output[6][19] , \stage_3_output[6][18] ,
         \stage_3_output[6][17] , \stage_3_output[6][16] ,
         \stage_3_output[6][15] , \stage_3_output[6][14] ,
         \stage_3_output[6][13] , \stage_3_output[6][12] ,
         \stage_3_output[6][11] , \stage_3_output[6][10] ,
         \stage_3_output[6][9] , \stage_3_output[6][8] ,
         \stage_3_output[6][7] , \stage_3_output[6][6] ,
         \stage_3_output[6][5] , \stage_3_output[6][4] ,
         \stage_3_output[6][3] , \stage_3_output[6][2] ,
         \stage_3_output[6][1] , \stage_3_output[6][0] ,
         \stage_3_output[5][19] , \stage_3_output[5][18] ,
         \stage_3_output[5][17] , \stage_3_output[5][16] ,
         \stage_3_output[5][15] , \stage_3_output[5][14] ,
         \stage_3_output[5][13] , \stage_3_output[5][12] ,
         \stage_3_output[5][11] , \stage_3_output[5][10] ,
         \stage_3_output[5][9] , \stage_3_output[5][8] ,
         \stage_3_output[5][7] , \stage_3_output[5][6] ,
         \stage_3_output[5][5] , \stage_3_output[5][4] ,
         \stage_3_output[5][3] , \stage_3_output[5][2] ,
         \stage_3_output[5][1] , \stage_3_output[5][0] ,
         \stage_3_output[4][19] , \stage_3_output[4][18] ,
         \stage_3_output[4][17] , \stage_3_output[4][16] ,
         \stage_3_output[4][15] , \stage_3_output[4][14] ,
         \stage_3_output[4][13] , \stage_3_output[4][12] ,
         \stage_3_output[4][11] , \stage_3_output[4][10] ,
         \stage_3_output[4][9] , \stage_3_output[4][8] ,
         \stage_3_output[4][7] , \stage_3_output[4][6] ,
         \stage_3_output[4][5] , \stage_3_output[4][4] ,
         \stage_3_output[4][3] , \stage_3_output[4][2] ,
         \stage_3_output[4][1] , \stage_3_output[4][0] ,
         \stage_3_output[3][19] , \stage_3_output[3][18] ,
         \stage_3_output[3][17] , \stage_3_output[3][16] ,
         \stage_3_output[3][15] , \stage_3_output[3][14] ,
         \stage_3_output[3][13] , \stage_3_output[3][12] ,
         \stage_3_output[3][11] , \stage_3_output[3][10] ,
         \stage_3_output[3][9] , \stage_3_output[3][8] ,
         \stage_3_output[3][7] , \stage_3_output[3][6] ,
         \stage_3_output[3][5] , \stage_3_output[3][4] ,
         \stage_3_output[3][3] , \stage_3_output[3][2] ,
         \stage_3_output[3][1] , \stage_3_output[3][0] ,
         \stage_3_output[2][19] , \stage_3_output[2][18] ,
         \stage_3_output[2][17] , \stage_3_output[2][16] ,
         \stage_3_output[2][15] , \stage_3_output[2][14] ,
         \stage_3_output[2][13] , \stage_3_output[2][12] ,
         \stage_3_output[2][11] , \stage_3_output[2][10] ,
         \stage_3_output[2][9] , \stage_3_output[2][8] ,
         \stage_3_output[2][7] , \stage_3_output[2][6] ,
         \stage_3_output[2][5] , \stage_3_output[2][4] ,
         \stage_3_output[2][3] , \stage_3_output[2][2] ,
         \stage_3_output[2][1] , \stage_3_output[2][0] ,
         \stage_3_output[1][19] , \stage_3_output[1][18] ,
         \stage_3_output[1][17] , \stage_3_output[1][16] ,
         \stage_3_output[1][15] , \stage_3_output[1][14] ,
         \stage_3_output[1][13] , \stage_3_output[1][12] ,
         \stage_3_output[1][11] , \stage_3_output[1][10] ,
         \stage_3_output[1][9] , \stage_3_output[1][8] ,
         \stage_3_output[1][7] , \stage_3_output[1][6] ,
         \stage_3_output[1][5] , \stage_3_output[1][4] ,
         \stage_3_output[1][3] , \stage_3_output[1][2] ,
         \stage_3_output[1][1] , \stage_3_output[1][0] ,
         \stage_3_output[0][19] , \stage_3_output[0][18] ,
         \stage_3_output[0][17] , \stage_3_output[0][16] ,
         \stage_3_output[0][15] , \stage_3_output[0][14] ,
         \stage_3_output[0][13] , \stage_3_output[0][12] ,
         \stage_3_output[0][11] , \stage_3_output[0][10] ,
         \stage_3_output[0][9] , \stage_3_output[0][8] ,
         \stage_3_output[0][7] , \stage_3_output[0][6] ,
         \stage_3_output[0][5] , \stage_3_output[0][4] ,
         \stage_3_output[0][3] , \stage_3_output[0][2] ,
         \stage_3_output[0][1] , \stage_3_output[0][0] ,
         \stage_3_retimer[7][19] , \stage_3_retimer[7][18] ,
         \stage_3_retimer[7][17] , \stage_3_retimer[7][16] ,
         \stage_3_retimer[7][15] , \stage_3_retimer[7][14] ,
         \stage_3_retimer[7][13] , \stage_3_retimer[7][12] ,
         \stage_3_retimer[7][11] , \stage_3_retimer[7][10] ,
         \stage_3_retimer[7][9] , \stage_3_retimer[7][8] ,
         \stage_3_retimer[7][7] , \stage_3_retimer[7][6] ,
         \stage_3_retimer[7][5] , \stage_3_retimer[7][4] ,
         \stage_3_retimer[7][3] , \stage_3_retimer[7][2] ,
         \stage_3_retimer[7][1] , \stage_3_retimer[7][0] ,
         \stage_3_retimer[6][19] , \stage_3_retimer[6][18] ,
         \stage_3_retimer[6][17] , \stage_3_retimer[6][16] ,
         \stage_3_retimer[6][15] , \stage_3_retimer[6][14] ,
         \stage_3_retimer[6][13] , \stage_3_retimer[6][12] ,
         \stage_3_retimer[6][11] , \stage_3_retimer[6][10] ,
         \stage_3_retimer[6][9] , \stage_3_retimer[6][8] ,
         \stage_3_retimer[6][7] , \stage_3_retimer[6][6] ,
         \stage_3_retimer[6][5] , \stage_3_retimer[6][4] ,
         \stage_3_retimer[6][3] , \stage_3_retimer[6][2] ,
         \stage_3_retimer[6][1] , \stage_3_retimer[6][0] ,
         \stage_3_retimer[5][19] , \stage_3_retimer[5][18] ,
         \stage_3_retimer[5][17] , \stage_3_retimer[5][16] ,
         \stage_3_retimer[5][15] , \stage_3_retimer[5][14] ,
         \stage_3_retimer[5][13] , \stage_3_retimer[5][12] ,
         \stage_3_retimer[5][11] , \stage_3_retimer[5][10] ,
         \stage_3_retimer[5][9] , \stage_3_retimer[5][8] ,
         \stage_3_retimer[5][7] , \stage_3_retimer[5][6] ,
         \stage_3_retimer[5][5] , \stage_3_retimer[5][4] ,
         \stage_3_retimer[5][3] , \stage_3_retimer[5][2] ,
         \stage_3_retimer[5][1] , \stage_3_retimer[5][0] ,
         \stage_3_retimer[4][19] , \stage_3_retimer[4][18] ,
         \stage_3_retimer[4][17] , \stage_3_retimer[4][16] ,
         \stage_3_retimer[4][15] , \stage_3_retimer[4][14] ,
         \stage_3_retimer[4][13] , \stage_3_retimer[4][12] ,
         \stage_3_retimer[4][11] , \stage_3_retimer[4][10] ,
         \stage_3_retimer[4][9] , \stage_3_retimer[4][8] ,
         \stage_3_retimer[4][7] , \stage_3_retimer[4][6] ,
         \stage_3_retimer[4][5] , \stage_3_retimer[4][4] ,
         \stage_3_retimer[4][3] , \stage_3_retimer[4][2] ,
         \stage_3_retimer[4][1] , \stage_3_retimer[4][0] ,
         \stage_3_retimer[3][19] , \stage_3_retimer[3][18] ,
         \stage_3_retimer[3][17] , \stage_3_retimer[3][16] ,
         \stage_3_retimer[3][15] , \stage_3_retimer[3][14] ,
         \stage_3_retimer[3][13] , \stage_3_retimer[3][12] ,
         \stage_3_retimer[3][11] , \stage_3_retimer[3][10] ,
         \stage_3_retimer[3][9] , \stage_3_retimer[3][8] ,
         \stage_3_retimer[3][7] , \stage_3_retimer[3][6] ,
         \stage_3_retimer[3][5] , \stage_3_retimer[3][4] ,
         \stage_3_retimer[3][3] , \stage_3_retimer[3][2] ,
         \stage_3_retimer[3][1] , \stage_3_retimer[3][0] ,
         \stage_3_retimer[2][19] , \stage_3_retimer[2][18] ,
         \stage_3_retimer[2][17] , \stage_3_retimer[2][16] ,
         \stage_3_retimer[2][15] , \stage_3_retimer[2][14] ,
         \stage_3_retimer[2][13] , \stage_3_retimer[2][12] ,
         \stage_3_retimer[2][11] , \stage_3_retimer[2][10] ,
         \stage_3_retimer[2][9] , \stage_3_retimer[2][8] ,
         \stage_3_retimer[2][7] , \stage_3_retimer[2][6] ,
         \stage_3_retimer[2][5] , \stage_3_retimer[2][4] ,
         \stage_3_retimer[2][3] , \stage_3_retimer[2][2] ,
         \stage_3_retimer[2][1] , \stage_3_retimer[2][0] ,
         \stage_3_retimer[1][19] , \stage_3_retimer[1][18] ,
         \stage_3_retimer[1][17] , \stage_3_retimer[1][16] ,
         \stage_3_retimer[1][15] , \stage_3_retimer[1][14] ,
         \stage_3_retimer[1][13] , \stage_3_retimer[1][12] ,
         \stage_3_retimer[1][11] , \stage_3_retimer[1][10] ,
         \stage_3_retimer[1][9] , \stage_3_retimer[1][8] ,
         \stage_3_retimer[1][7] , \stage_3_retimer[1][6] ,
         \stage_3_retimer[1][5] , \stage_3_retimer[1][4] ,
         \stage_3_retimer[1][3] , \stage_3_retimer[1][2] ,
         \stage_3_retimer[1][1] , \stage_3_retimer[1][0] ,
         \stage_3_retimer[0][19] , \stage_3_retimer[0][18] ,
         \stage_3_retimer[0][17] , \stage_3_retimer[0][16] ,
         \stage_3_retimer[0][15] , \stage_3_retimer[0][14] ,
         \stage_3_retimer[0][13] , \stage_3_retimer[0][12] ,
         \stage_3_retimer[0][11] , \stage_3_retimer[0][10] ,
         \stage_3_retimer[0][9] , \stage_3_retimer[0][8] ,
         \stage_3_retimer[0][7] , \stage_3_retimer[0][6] ,
         \stage_3_retimer[0][5] , \stage_3_retimer[0][4] ,
         \stage_3_retimer[0][3] , \stage_3_retimer[0][2] ,
         \stage_3_retimer[0][1] , \stage_3_retimer[0][0] ,
         \stage_4_output[7][19] , \stage_4_output[7][18] ,
         \stage_4_output[7][17] , \stage_4_output[7][16] ,
         \stage_4_output[7][15] , \stage_4_output[7][14] ,
         \stage_4_output[7][13] , \stage_4_output[7][12] ,
         \stage_4_output[7][11] , \stage_4_output[7][10] ,
         \stage_4_output[7][9] , \stage_4_output[7][8] ,
         \stage_4_output[7][7] , \stage_4_output[7][6] ,
         \stage_4_output[7][5] , \stage_4_output[7][4] ,
         \stage_4_output[7][3] , \stage_4_output[7][2] ,
         \stage_4_output[7][1] , \stage_4_output[7][0] ,
         \stage_4_output[6][19] , \stage_4_output[6][18] ,
         \stage_4_output[6][17] , \stage_4_output[6][16] ,
         \stage_4_output[6][15] , \stage_4_output[6][14] ,
         \stage_4_output[6][13] , \stage_4_output[6][12] ,
         \stage_4_output[6][11] , \stage_4_output[6][10] ,
         \stage_4_output[6][9] , \stage_4_output[6][8] ,
         \stage_4_output[6][7] , \stage_4_output[6][6] ,
         \stage_4_output[6][5] , \stage_4_output[6][4] ,
         \stage_4_output[6][3] , \stage_4_output[6][2] ,
         \stage_4_output[6][1] , \stage_4_output[6][0] ,
         \stage_4_output[5][19] , \stage_4_output[5][18] ,
         \stage_4_output[5][17] , \stage_4_output[5][16] ,
         \stage_4_output[5][15] , \stage_4_output[5][14] ,
         \stage_4_output[5][13] , \stage_4_output[5][12] ,
         \stage_4_output[5][11] , \stage_4_output[5][10] ,
         \stage_4_output[5][9] , \stage_4_output[5][8] ,
         \stage_4_output[5][7] , \stage_4_output[5][6] ,
         \stage_4_output[5][5] , \stage_4_output[5][4] ,
         \stage_4_output[5][3] , \stage_4_output[5][2] ,
         \stage_4_output[5][1] , \stage_4_output[5][0] ,
         \stage_4_output[4][19] , \stage_4_output[4][18] ,
         \stage_4_output[4][17] , \stage_4_output[4][16] ,
         \stage_4_output[4][15] , \stage_4_output[4][14] ,
         \stage_4_output[4][13] , \stage_4_output[4][12] ,
         \stage_4_output[4][11] , \stage_4_output[4][10] ,
         \stage_4_output[4][9] , \stage_4_output[4][8] ,
         \stage_4_output[4][7] , \stage_4_output[4][6] ,
         \stage_4_output[4][5] , \stage_4_output[4][4] ,
         \stage_4_output[4][3] , \stage_4_output[4][2] ,
         \stage_4_output[4][1] , \stage_4_output[4][0] ,
         \stage_4_output[3][19] , \stage_4_output[3][18] ,
         \stage_4_output[3][17] , \stage_4_output[3][16] ,
         \stage_4_output[3][15] , \stage_4_output[3][14] ,
         \stage_4_output[3][13] , \stage_4_output[3][12] ,
         \stage_4_output[3][11] , \stage_4_output[3][10] ,
         \stage_4_output[3][9] , \stage_4_output[3][8] ,
         \stage_4_output[3][7] , \stage_4_output[3][6] ,
         \stage_4_output[3][5] , \stage_4_output[3][4] ,
         \stage_4_output[3][3] , \stage_4_output[3][2] ,
         \stage_4_output[3][1] , \stage_4_output[3][0] ,
         \stage_4_output[2][19] , \stage_4_output[2][18] ,
         \stage_4_output[2][17] , \stage_4_output[2][16] ,
         \stage_4_output[2][15] , \stage_4_output[2][14] ,
         \stage_4_output[2][13] , \stage_4_output[2][12] ,
         \stage_4_output[2][11] , \stage_4_output[2][10] ,
         \stage_4_output[2][9] , \stage_4_output[2][8] ,
         \stage_4_output[2][7] , \stage_4_output[2][6] ,
         \stage_4_output[2][5] , \stage_4_output[2][4] ,
         \stage_4_output[2][3] , \stage_4_output[2][2] ,
         \stage_4_output[2][1] , \stage_4_output[2][0] ,
         \stage_4_output[1][19] , \stage_4_output[1][18] ,
         \stage_4_output[1][17] , \stage_4_output[1][16] ,
         \stage_4_output[1][15] , \stage_4_output[1][14] ,
         \stage_4_output[1][13] , \stage_4_output[1][12] ,
         \stage_4_output[1][11] , \stage_4_output[1][10] ,
         \stage_4_output[1][9] , \stage_4_output[1][8] ,
         \stage_4_output[1][7] , \stage_4_output[1][6] ,
         \stage_4_output[1][5] , \stage_4_output[1][4] ,
         \stage_4_output[1][3] , \stage_4_output[1][2] ,
         \stage_4_output[1][1] , \stage_4_output[1][0] ,
         \stage_4_output[0][19] , \stage_4_output[0][18] ,
         \stage_4_output[0][17] , \stage_4_output[0][16] ,
         \stage_4_output[0][15] , \stage_4_output[0][14] ,
         \stage_4_output[0][13] , \stage_4_output[0][12] ,
         \stage_4_output[0][11] , \stage_4_output[0][10] ,
         \stage_4_output[0][9] , \stage_4_output[0][8] ,
         \stage_4_output[0][7] , \stage_4_output[0][6] ,
         \stage_4_output[0][5] , \stage_4_output[0][4] ,
         \stage_4_output[0][3] , \stage_4_output[0][2] ,
         \stage_4_output[0][1] , \stage_4_output[0][0] ;
  assign \in_upper_00[3]  = port_en_n[0];
  assign \in_lower_00[3]  = port_en_n[1];
  assign \in_upper_01[3]  = port_en_n[2];
  assign \in_lower_01[3]  = port_en_n[3];
  assign in_upper_02_3 = port_en_n[4];
  assign \in_lower_02[3]  = port_en_n[5];
  assign \in_upper_03[3]  = port_en_n[6];

  crossbar_0 u_00_crossbar ( .in_upper({in_input[127:112], \in_upper_00[3] , 
        \in_upper_00[3] , \in_upper_00[3] , \in_upper_00[3] }), .in_lower({
        in_input[111:96], \in_lower_00[3] , \in_lower_00[3] , \in_lower_00[3] , 
        \*Logic1* }), .in_control(in_control[19]), .out_upper({
        \stage_0_output[0][19] , \stage_0_output[0][18] , 
        \stage_0_output[0][17] , \stage_0_output[0][16] , 
        \stage_0_output[0][15] , \stage_0_output[0][14] , 
        \stage_0_output[0][13] , \stage_0_output[0][12] , 
        \stage_0_output[0][11] , \stage_0_output[0][10] , 
        \stage_0_output[0][9] , \stage_0_output[0][8] , \stage_0_output[0][7] , 
        \stage_0_output[0][6] , \stage_0_output[0][5] , \stage_0_output[0][4] , 
        \stage_0_output[0][3] , \stage_0_output[0][2] , \stage_0_output[0][1] , 
        \stage_0_output[0][0] }), .out_lower({\stage_0_output[1][19] , 
        \stage_0_output[1][18] , \stage_0_output[1][17] , 
        \stage_0_output[1][16] , \stage_0_output[1][15] , 
        \stage_0_output[1][14] , \stage_0_output[1][13] , 
        \stage_0_output[1][12] , \stage_0_output[1][11] , 
        \stage_0_output[1][10] , \stage_0_output[1][9] , 
        \stage_0_output[1][8] , \stage_0_output[1][7] , \stage_0_output[1][6] , 
        \stage_0_output[1][5] , \stage_0_output[1][4] , \stage_0_output[1][3] , 
        \stage_0_output[1][2] , \stage_0_output[1][1] , \stage_0_output[1][0] }) );
  crossbar_19 u_01_crossbar ( .in_upper({in_input[95:80], \in_upper_01[3] , 
        \in_upper_01[3] , \*Logic1* , \in_upper_01[3] }), .in_lower({
        in_input[79:64], \in_lower_01[3] , \in_lower_01[3] , \*Logic1* , 
        \*Logic1* }), .in_control(in_control[18]), .out_upper({
        \stage_0_output[2][19] , \stage_0_output[2][18] , 
        \stage_0_output[2][17] , \stage_0_output[2][16] , 
        \stage_0_output[2][15] , \stage_0_output[2][14] , 
        \stage_0_output[2][13] , \stage_0_output[2][12] , 
        \stage_0_output[2][11] , \stage_0_output[2][10] , 
        \stage_0_output[2][9] , \stage_0_output[2][8] , \stage_0_output[2][7] , 
        \stage_0_output[2][6] , \stage_0_output[2][5] , \stage_0_output[2][4] , 
        \stage_0_output[2][3] , \stage_0_output[2][2] , \stage_0_output[2][1] , 
        \stage_0_output[2][0] }), .out_lower({\stage_0_output[3][19] , 
        \stage_0_output[3][18] , \stage_0_output[3][17] , 
        \stage_0_output[3][16] , \stage_0_output[3][15] , 
        \stage_0_output[3][14] , \stage_0_output[3][13] , 
        \stage_0_output[3][12] , \stage_0_output[3][11] , 
        \stage_0_output[3][10] , \stage_0_output[3][9] , 
        \stage_0_output[3][8] , \stage_0_output[3][7] , \stage_0_output[3][6] , 
        \stage_0_output[3][5] , \stage_0_output[3][4] , \stage_0_output[3][3] , 
        \stage_0_output[3][2] , \stage_0_output[3][1] , \stage_0_output[3][0] }) );
  crossbar_18 u_02_crossbar ( .in_upper({in_input[63:48], in_upper_02_3, 
        \*Logic1* , in_upper_02_3, in_upper_02_3}), .in_lower({in_input[47:32], 
        \in_lower_02[3] , \*Logic1* , \in_lower_02[3] , \*Logic1* }), 
        .in_control(in_control[17]), .out_upper({\stage_0_output[4][19] , 
        \stage_0_output[4][18] , \stage_0_output[4][17] , 
        \stage_0_output[4][16] , \stage_0_output[4][15] , 
        \stage_0_output[4][14] , \stage_0_output[4][13] , 
        \stage_0_output[4][12] , \stage_0_output[4][11] , 
        \stage_0_output[4][10] , \stage_0_output[4][9] , 
        \stage_0_output[4][8] , \stage_0_output[4][7] , \stage_0_output[4][6] , 
        \stage_0_output[4][5] , \stage_0_output[4][4] , \stage_0_output[4][3] , 
        \stage_0_output[4][2] , \stage_0_output[4][1] , \stage_0_output[4][0] }), .out_lower({\stage_0_output[5][19] , \stage_0_output[5][18] , 
        \stage_0_output[5][17] , \stage_0_output[5][16] , 
        \stage_0_output[5][15] , \stage_0_output[5][14] , 
        \stage_0_output[5][13] , \stage_0_output[5][12] , 
        \stage_0_output[5][11] , \stage_0_output[5][10] , 
        \stage_0_output[5][9] , \stage_0_output[5][8] , \stage_0_output[5][7] , 
        \stage_0_output[5][6] , \stage_0_output[5][5] , \stage_0_output[5][4] , 
        \stage_0_output[5][3] , \stage_0_output[5][2] , \stage_0_output[5][1] , 
        \stage_0_output[5][0] }) );
  crossbar_17 u_03_crossbar ( .in_upper({in_input[31:16], \in_upper_03[3] , 
        \*Logic1* , \*Logic1* , \in_upper_03[3] }), .in_lower({in_input[15:0], 
        port_en_n[7], \*Logic1* , \*Logic1* , \*Logic1* }), .in_control(
        in_control[16]), .out_upper({\stage_0_output[6][19] , 
        \stage_0_output[6][18] , \stage_0_output[6][17] , 
        \stage_0_output[6][16] , \stage_0_output[6][15] , 
        \stage_0_output[6][14] , \stage_0_output[6][13] , 
        \stage_0_output[6][12] , \stage_0_output[6][11] , 
        \stage_0_output[6][10] , \stage_0_output[6][9] , 
        \stage_0_output[6][8] , \stage_0_output[6][7] , \stage_0_output[6][6] , 
        \stage_0_output[6][5] , \stage_0_output[6][4] , \stage_0_output[6][3] , 
        \stage_0_output[6][2] , \stage_0_output[6][1] , \stage_0_output[6][0] }), .out_lower({\stage_0_output[7][19] , \stage_0_output[7][18] , 
        \stage_0_output[7][17] , \stage_0_output[7][16] , 
        \stage_0_output[7][15] , \stage_0_output[7][14] , 
        \stage_0_output[7][13] , \stage_0_output[7][12] , 
        \stage_0_output[7][11] , \stage_0_output[7][10] , 
        \stage_0_output[7][9] , \stage_0_output[7][8] , \stage_0_output[7][7] , 
        \stage_0_output[7][6] , \stage_0_output[7][5] , \stage_0_output[7][4] , 
        \stage_0_output[7][3] , \stage_0_output[7][2] , \stage_0_output[7][1] , 
        \stage_0_output[7][0] }) );
  crossbar_16 u_10_crossbar ( .in_upper({\stage_0_retimer[0][19] , 
        \stage_0_retimer[0][18] , \stage_0_retimer[0][17] , 
        \stage_0_retimer[0][16] , \stage_0_retimer[0][15] , 
        \stage_0_retimer[0][14] , \stage_0_retimer[0][13] , 
        \stage_0_retimer[0][12] , \stage_0_retimer[0][11] , 
        \stage_0_retimer[0][10] , \stage_0_retimer[0][9] , 
        \stage_0_retimer[0][8] , \stage_0_retimer[0][7] , 
        \stage_0_retimer[0][6] , \stage_0_retimer[0][5] , 
        \stage_0_retimer[0][4] , \stage_0_retimer[0][3] , 
        \stage_0_retimer[0][2] , \stage_0_retimer[0][1] , 
        \stage_0_retimer[0][0] }), .in_lower({\stage_0_retimer[2][19] , 
        \stage_0_retimer[2][18] , \stage_0_retimer[2][17] , 
        \stage_0_retimer[2][16] , \stage_0_retimer[2][15] , 
        \stage_0_retimer[2][14] , \stage_0_retimer[2][13] , 
        \stage_0_retimer[2][12] , \stage_0_retimer[2][11] , 
        \stage_0_retimer[2][10] , \stage_0_retimer[2][9] , 
        \stage_0_retimer[2][8] , \stage_0_retimer[2][7] , 
        \stage_0_retimer[2][6] , \stage_0_retimer[2][5] , 
        \stage_0_retimer[2][4] , \stage_0_retimer[2][3] , 
        \stage_0_retimer[2][2] , \stage_0_retimer[2][1] , 
        \stage_0_retimer[2][0] }), .in_control(in_control[15]), .out_upper({
        \stage_1_output[0][19] , \stage_1_output[0][18] , 
        \stage_1_output[0][17] , \stage_1_output[0][16] , 
        \stage_1_output[0][15] , \stage_1_output[0][14] , 
        \stage_1_output[0][13] , \stage_1_output[0][12] , 
        \stage_1_output[0][11] , \stage_1_output[0][10] , 
        \stage_1_output[0][9] , \stage_1_output[0][8] , \stage_1_output[0][7] , 
        \stage_1_output[0][6] , \stage_1_output[0][5] , \stage_1_output[0][4] , 
        \stage_1_output[0][3] , \stage_1_output[0][2] , \stage_1_output[0][1] , 
        \stage_1_output[0][0] }), .out_lower({\stage_1_output[1][19] , 
        \stage_1_output[1][18] , \stage_1_output[1][17] , 
        \stage_1_output[1][16] , \stage_1_output[1][15] , 
        \stage_1_output[1][14] , \stage_1_output[1][13] , 
        \stage_1_output[1][12] , \stage_1_output[1][11] , 
        \stage_1_output[1][10] , \stage_1_output[1][9] , 
        \stage_1_output[1][8] , \stage_1_output[1][7] , \stage_1_output[1][6] , 
        \stage_1_output[1][5] , \stage_1_output[1][4] , \stage_1_output[1][3] , 
        \stage_1_output[1][2] , \stage_1_output[1][1] , \stage_1_output[1][0] }) );
  crossbar_15 u_11_crossbar ( .in_upper({\stage_0_retimer[4][19] , 
        \stage_0_retimer[4][18] , \stage_0_retimer[4][17] , 
        \stage_0_retimer[4][16] , \stage_0_retimer[4][15] , 
        \stage_0_retimer[4][14] , \stage_0_retimer[4][13] , 
        \stage_0_retimer[4][12] , \stage_0_retimer[4][11] , 
        \stage_0_retimer[4][10] , \stage_0_retimer[4][9] , 
        \stage_0_retimer[4][8] , \stage_0_retimer[4][7] , 
        \stage_0_retimer[4][6] , \stage_0_retimer[4][5] , 
        \stage_0_retimer[4][4] , \stage_0_retimer[4][3] , 
        \stage_0_retimer[4][2] , \stage_0_retimer[4][1] , 
        \stage_0_retimer[4][0] }), .in_lower({\stage_0_retimer[6][19] , 
        \stage_0_retimer[6][18] , \stage_0_retimer[6][17] , 
        \stage_0_retimer[6][16] , \stage_0_retimer[6][15] , 
        \stage_0_retimer[6][14] , \stage_0_retimer[6][13] , 
        \stage_0_retimer[6][12] , \stage_0_retimer[6][11] , 
        \stage_0_retimer[6][10] , \stage_0_retimer[6][9] , 
        \stage_0_retimer[6][8] , \stage_0_retimer[6][7] , 
        \stage_0_retimer[6][6] , \stage_0_retimer[6][5] , 
        \stage_0_retimer[6][4] , \stage_0_retimer[6][3] , 
        \stage_0_retimer[6][2] , \stage_0_retimer[6][1] , 
        \stage_0_retimer[6][0] }), .in_control(in_control[14]), .out_upper({
        \stage_1_output[2][19] , \stage_1_output[2][18] , 
        \stage_1_output[2][17] , \stage_1_output[2][16] , 
        \stage_1_output[2][15] , \stage_1_output[2][14] , 
        \stage_1_output[2][13] , \stage_1_output[2][12] , 
        \stage_1_output[2][11] , \stage_1_output[2][10] , 
        \stage_1_output[2][9] , \stage_1_output[2][8] , \stage_1_output[2][7] , 
        \stage_1_output[2][6] , \stage_1_output[2][5] , \stage_1_output[2][4] , 
        \stage_1_output[2][3] , \stage_1_output[2][2] , \stage_1_output[2][1] , 
        \stage_1_output[2][0] }), .out_lower({\stage_1_output[3][19] , 
        \stage_1_output[3][18] , \stage_1_output[3][17] , 
        \stage_1_output[3][16] , \stage_1_output[3][15] , 
        \stage_1_output[3][14] , \stage_1_output[3][13] , 
        \stage_1_output[3][12] , \stage_1_output[3][11] , 
        \stage_1_output[3][10] , \stage_1_output[3][9] , 
        \stage_1_output[3][8] , \stage_1_output[3][7] , \stage_1_output[3][6] , 
        \stage_1_output[3][5] , \stage_1_output[3][4] , \stage_1_output[3][3] , 
        \stage_1_output[3][2] , \stage_1_output[3][1] , \stage_1_output[3][0] }) );
  crossbar_14 u_12_crossbar ( .in_upper({\stage_0_retimer[1][19] , 
        \stage_0_retimer[1][18] , \stage_0_retimer[1][17] , 
        \stage_0_retimer[1][16] , \stage_0_retimer[1][15] , 
        \stage_0_retimer[1][14] , \stage_0_retimer[1][13] , 
        \stage_0_retimer[1][12] , \stage_0_retimer[1][11] , 
        \stage_0_retimer[1][10] , \stage_0_retimer[1][9] , 
        \stage_0_retimer[1][8] , \stage_0_retimer[1][7] , 
        \stage_0_retimer[1][6] , \stage_0_retimer[1][5] , 
        \stage_0_retimer[1][4] , \stage_0_retimer[1][3] , 
        \stage_0_retimer[1][2] , \stage_0_retimer[1][1] , 
        \stage_0_retimer[1][0] }), .in_lower({\stage_0_retimer[3][19] , 
        \stage_0_retimer[3][18] , \stage_0_retimer[3][17] , 
        \stage_0_retimer[3][16] , \stage_0_retimer[3][15] , 
        \stage_0_retimer[3][14] , \stage_0_retimer[3][13] , 
        \stage_0_retimer[3][12] , \stage_0_retimer[3][11] , 
        \stage_0_retimer[3][10] , \stage_0_retimer[3][9] , 
        \stage_0_retimer[3][8] , \stage_0_retimer[3][7] , 
        \stage_0_retimer[3][6] , \stage_0_retimer[3][5] , 
        \stage_0_retimer[3][4] , \stage_0_retimer[3][3] , 
        \stage_0_retimer[3][2] , \stage_0_retimer[3][1] , 
        \stage_0_retimer[3][0] }), .in_control(in_control[13]), .out_upper({
        \stage_1_output[4][19] , \stage_1_output[4][18] , 
        \stage_1_output[4][17] , \stage_1_output[4][16] , 
        \stage_1_output[4][15] , \stage_1_output[4][14] , 
        \stage_1_output[4][13] , \stage_1_output[4][12] , 
        \stage_1_output[4][11] , \stage_1_output[4][10] , 
        \stage_1_output[4][9] , \stage_1_output[4][8] , \stage_1_output[4][7] , 
        \stage_1_output[4][6] , \stage_1_output[4][5] , \stage_1_output[4][4] , 
        \stage_1_output[4][3] , \stage_1_output[4][2] , \stage_1_output[4][1] , 
        \stage_1_output[4][0] }), .out_lower({\stage_1_output[5][19] , 
        \stage_1_output[5][18] , \stage_1_output[5][17] , 
        \stage_1_output[5][16] , \stage_1_output[5][15] , 
        \stage_1_output[5][14] , \stage_1_output[5][13] , 
        \stage_1_output[5][12] , \stage_1_output[5][11] , 
        \stage_1_output[5][10] , \stage_1_output[5][9] , 
        \stage_1_output[5][8] , \stage_1_output[5][7] , \stage_1_output[5][6] , 
        \stage_1_output[5][5] , \stage_1_output[5][4] , \stage_1_output[5][3] , 
        \stage_1_output[5][2] , \stage_1_output[5][1] , \stage_1_output[5][0] }) );
  crossbar_13 u_13_crossbar ( .in_upper({\stage_0_retimer[5][19] , 
        \stage_0_retimer[5][18] , \stage_0_retimer[5][17] , 
        \stage_0_retimer[5][16] , \stage_0_retimer[5][15] , 
        \stage_0_retimer[5][14] , \stage_0_retimer[5][13] , 
        \stage_0_retimer[5][12] , \stage_0_retimer[5][11] , 
        \stage_0_retimer[5][10] , \stage_0_retimer[5][9] , 
        \stage_0_retimer[5][8] , \stage_0_retimer[5][7] , 
        \stage_0_retimer[5][6] , \stage_0_retimer[5][5] , 
        \stage_0_retimer[5][4] , \stage_0_retimer[5][3] , 
        \stage_0_retimer[5][2] , \stage_0_retimer[5][1] , 
        \stage_0_retimer[5][0] }), .in_lower({\stage_0_retimer[7][19] , 
        \stage_0_retimer[7][18] , \stage_0_retimer[7][17] , 
        \stage_0_retimer[7][16] , \stage_0_retimer[7][15] , 
        \stage_0_retimer[7][14] , \stage_0_retimer[7][13] , 
        \stage_0_retimer[7][12] , \stage_0_retimer[7][11] , 
        \stage_0_retimer[7][10] , \stage_0_retimer[7][9] , 
        \stage_0_retimer[7][8] , \stage_0_retimer[7][7] , 
        \stage_0_retimer[7][6] , \stage_0_retimer[7][5] , 
        \stage_0_retimer[7][4] , \stage_0_retimer[7][3] , 
        \stage_0_retimer[7][2] , \stage_0_retimer[7][1] , 
        \stage_0_retimer[7][0] }), .in_control(in_control[12]), .out_upper({
        \stage_1_output[6][19] , \stage_1_output[6][18] , 
        \stage_1_output[6][17] , \stage_1_output[6][16] , 
        \stage_1_output[6][15] , \stage_1_output[6][14] , 
        \stage_1_output[6][13] , \stage_1_output[6][12] , 
        \stage_1_output[6][11] , \stage_1_output[6][10] , 
        \stage_1_output[6][9] , \stage_1_output[6][8] , \stage_1_output[6][7] , 
        \stage_1_output[6][6] , \stage_1_output[6][5] , \stage_1_output[6][4] , 
        \stage_1_output[6][3] , \stage_1_output[6][2] , \stage_1_output[6][1] , 
        \stage_1_output[6][0] }), .out_lower({\stage_1_output[7][19] , 
        \stage_1_output[7][18] , \stage_1_output[7][17] , 
        \stage_1_output[7][16] , \stage_1_output[7][15] , 
        \stage_1_output[7][14] , \stage_1_output[7][13] , 
        \stage_1_output[7][12] , \stage_1_output[7][11] , 
        \stage_1_output[7][10] , \stage_1_output[7][9] , 
        \stage_1_output[7][8] , \stage_1_output[7][7] , \stage_1_output[7][6] , 
        \stage_1_output[7][5] , \stage_1_output[7][4] , \stage_1_output[7][3] , 
        \stage_1_output[7][2] , \stage_1_output[7][1] , \stage_1_output[7][0] }) );
  crossbar_12 u_20_crossbar ( .in_upper({\stage_1_retimer[0][19] , 
        \stage_1_retimer[0][18] , \stage_1_retimer[0][17] , 
        \stage_1_retimer[0][16] , \stage_1_retimer[0][15] , 
        \stage_1_retimer[0][14] , \stage_1_retimer[0][13] , 
        \stage_1_retimer[0][12] , \stage_1_retimer[0][11] , 
        \stage_1_retimer[0][10] , \stage_1_retimer[0][9] , 
        \stage_1_retimer[0][8] , \stage_1_retimer[0][7] , 
        \stage_1_retimer[0][6] , \stage_1_retimer[0][5] , 
        \stage_1_retimer[0][4] , \stage_1_retimer[0][3] , 
        \stage_1_retimer[0][2] , \stage_1_retimer[0][1] , 
        \stage_1_retimer[0][0] }), .in_lower({\stage_1_retimer[2][19] , 
        \stage_1_retimer[2][18] , \stage_1_retimer[2][17] , 
        \stage_1_retimer[2][16] , \stage_1_retimer[2][15] , 
        \stage_1_retimer[2][14] , \stage_1_retimer[2][13] , 
        \stage_1_retimer[2][12] , \stage_1_retimer[2][11] , 
        \stage_1_retimer[2][10] , \stage_1_retimer[2][9] , 
        \stage_1_retimer[2][8] , \stage_1_retimer[2][7] , 
        \stage_1_retimer[2][6] , \stage_1_retimer[2][5] , 
        \stage_1_retimer[2][4] , \stage_1_retimer[2][3] , 
        \stage_1_retimer[2][2] , \stage_1_retimer[2][1] , 
        \stage_1_retimer[2][0] }), .in_control(in_control[11]), .out_upper({
        \stage_2_output[0][19] , \stage_2_output[0][18] , 
        \stage_2_output[0][17] , \stage_2_output[0][16] , 
        \stage_2_output[0][15] , \stage_2_output[0][14] , 
        \stage_2_output[0][13] , \stage_2_output[0][12] , 
        \stage_2_output[0][11] , \stage_2_output[0][10] , 
        \stage_2_output[0][9] , \stage_2_output[0][8] , \stage_2_output[0][7] , 
        \stage_2_output[0][6] , \stage_2_output[0][5] , \stage_2_output[0][4] , 
        \stage_2_output[0][3] , \stage_2_output[0][2] , \stage_2_output[0][1] , 
        \stage_2_output[0][0] }), .out_lower({\stage_2_output[1][19] , 
        \stage_2_output[1][18] , \stage_2_output[1][17] , 
        \stage_2_output[1][16] , \stage_2_output[1][15] , 
        \stage_2_output[1][14] , \stage_2_output[1][13] , 
        \stage_2_output[1][12] , \stage_2_output[1][11] , 
        \stage_2_output[1][10] , \stage_2_output[1][9] , 
        \stage_2_output[1][8] , \stage_2_output[1][7] , \stage_2_output[1][6] , 
        \stage_2_output[1][5] , \stage_2_output[1][4] , \stage_2_output[1][3] , 
        \stage_2_output[1][2] , \stage_2_output[1][1] , \stage_2_output[1][0] }) );
  crossbar_11 u_21_crossbar ( .in_upper({\stage_1_retimer[1][19] , 
        \stage_1_retimer[1][18] , \stage_1_retimer[1][17] , 
        \stage_1_retimer[1][16] , \stage_1_retimer[1][15] , 
        \stage_1_retimer[1][14] , \stage_1_retimer[1][13] , 
        \stage_1_retimer[1][12] , \stage_1_retimer[1][11] , 
        \stage_1_retimer[1][10] , \stage_1_retimer[1][9] , 
        \stage_1_retimer[1][8] , \stage_1_retimer[1][7] , 
        \stage_1_retimer[1][6] , \stage_1_retimer[1][5] , 
        \stage_1_retimer[1][4] , \stage_1_retimer[1][3] , 
        \stage_1_retimer[1][2] , \stage_1_retimer[1][1] , 
        \stage_1_retimer[1][0] }), .in_lower({\stage_1_retimer[3][19] , 
        \stage_1_retimer[3][18] , \stage_1_retimer[3][17] , 
        \stage_1_retimer[3][16] , \stage_1_retimer[3][15] , 
        \stage_1_retimer[3][14] , \stage_1_retimer[3][13] , 
        \stage_1_retimer[3][12] , \stage_1_retimer[3][11] , 
        \stage_1_retimer[3][10] , \stage_1_retimer[3][9] , 
        \stage_1_retimer[3][8] , \stage_1_retimer[3][7] , 
        \stage_1_retimer[3][6] , \stage_1_retimer[3][5] , 
        \stage_1_retimer[3][4] , \stage_1_retimer[3][3] , 
        \stage_1_retimer[3][2] , \stage_1_retimer[3][1] , 
        \stage_1_retimer[3][0] }), .in_control(in_control[10]), .out_upper({
        \stage_2_output[2][19] , \stage_2_output[2][18] , 
        \stage_2_output[2][17] , \stage_2_output[2][16] , 
        \stage_2_output[2][15] , \stage_2_output[2][14] , 
        \stage_2_output[2][13] , \stage_2_output[2][12] , 
        \stage_2_output[2][11] , \stage_2_output[2][10] , 
        \stage_2_output[2][9] , \stage_2_output[2][8] , \stage_2_output[2][7] , 
        \stage_2_output[2][6] , \stage_2_output[2][5] , \stage_2_output[2][4] , 
        \stage_2_output[2][3] , \stage_2_output[2][2] , \stage_2_output[2][1] , 
        \stage_2_output[2][0] }), .out_lower({\stage_2_output[3][19] , 
        \stage_2_output[3][18] , \stage_2_output[3][17] , 
        \stage_2_output[3][16] , \stage_2_output[3][15] , 
        \stage_2_output[3][14] , \stage_2_output[3][13] , 
        \stage_2_output[3][12] , \stage_2_output[3][11] , 
        \stage_2_output[3][10] , \stage_2_output[3][9] , 
        \stage_2_output[3][8] , \stage_2_output[3][7] , \stage_2_output[3][6] , 
        \stage_2_output[3][5] , \stage_2_output[3][4] , \stage_2_output[3][3] , 
        \stage_2_output[3][2] , \stage_2_output[3][1] , \stage_2_output[3][0] }) );
  crossbar_10 u_22_crossbar ( .in_upper({\stage_1_retimer[4][19] , 
        \stage_1_retimer[4][18] , \stage_1_retimer[4][17] , 
        \stage_1_retimer[4][16] , \stage_1_retimer[4][15] , 
        \stage_1_retimer[4][14] , \stage_1_retimer[4][13] , 
        \stage_1_retimer[4][12] , \stage_1_retimer[4][11] , 
        \stage_1_retimer[4][10] , \stage_1_retimer[4][9] , 
        \stage_1_retimer[4][8] , \stage_1_retimer[4][7] , 
        \stage_1_retimer[4][6] , \stage_1_retimer[4][5] , 
        \stage_1_retimer[4][4] , \stage_1_retimer[4][3] , 
        \stage_1_retimer[4][2] , \stage_1_retimer[4][1] , 
        \stage_1_retimer[4][0] }), .in_lower({\stage_1_retimer[6][19] , 
        \stage_1_retimer[6][18] , \stage_1_retimer[6][17] , 
        \stage_1_retimer[6][16] , \stage_1_retimer[6][15] , 
        \stage_1_retimer[6][14] , \stage_1_retimer[6][13] , 
        \stage_1_retimer[6][12] , \stage_1_retimer[6][11] , 
        \stage_1_retimer[6][10] , \stage_1_retimer[6][9] , 
        \stage_1_retimer[6][8] , \stage_1_retimer[6][7] , 
        \stage_1_retimer[6][6] , \stage_1_retimer[6][5] , 
        \stage_1_retimer[6][4] , \stage_1_retimer[6][3] , 
        \stage_1_retimer[6][2] , \stage_1_retimer[6][1] , 
        \stage_1_retimer[6][0] }), .in_control(in_control[9]), .out_upper({
        \stage_2_output[4][19] , \stage_2_output[4][18] , 
        \stage_2_output[4][17] , \stage_2_output[4][16] , 
        \stage_2_output[4][15] , \stage_2_output[4][14] , 
        \stage_2_output[4][13] , \stage_2_output[4][12] , 
        \stage_2_output[4][11] , \stage_2_output[4][10] , 
        \stage_2_output[4][9] , \stage_2_output[4][8] , \stage_2_output[4][7] , 
        \stage_2_output[4][6] , \stage_2_output[4][5] , \stage_2_output[4][4] , 
        \stage_2_output[4][3] , \stage_2_output[4][2] , \stage_2_output[4][1] , 
        \stage_2_output[4][0] }), .out_lower({\stage_2_output[5][19] , 
        \stage_2_output[5][18] , \stage_2_output[5][17] , 
        \stage_2_output[5][16] , \stage_2_output[5][15] , 
        \stage_2_output[5][14] , \stage_2_output[5][13] , 
        \stage_2_output[5][12] , \stage_2_output[5][11] , 
        \stage_2_output[5][10] , \stage_2_output[5][9] , 
        \stage_2_output[5][8] , \stage_2_output[5][7] , \stage_2_output[5][6] , 
        \stage_2_output[5][5] , \stage_2_output[5][4] , \stage_2_output[5][3] , 
        \stage_2_output[5][2] , \stage_2_output[5][1] , \stage_2_output[5][0] }) );
  crossbar_9 u_23_crossbar ( .in_upper({\stage_1_retimer[5][19] , 
        \stage_1_retimer[5][18] , \stage_1_retimer[5][17] , 
        \stage_1_retimer[5][16] , \stage_1_retimer[5][15] , 
        \stage_1_retimer[5][14] , \stage_1_retimer[5][13] , 
        \stage_1_retimer[5][12] , \stage_1_retimer[5][11] , 
        \stage_1_retimer[5][10] , \stage_1_retimer[5][9] , 
        \stage_1_retimer[5][8] , \stage_1_retimer[5][7] , 
        \stage_1_retimer[5][6] , \stage_1_retimer[5][5] , 
        \stage_1_retimer[5][4] , \stage_1_retimer[5][3] , 
        \stage_1_retimer[5][2] , \stage_1_retimer[5][1] , 
        \stage_1_retimer[5][0] }), .in_lower({\stage_1_retimer[7][19] , 
        \stage_1_retimer[7][18] , \stage_1_retimer[7][17] , 
        \stage_1_retimer[7][16] , \stage_1_retimer[7][15] , 
        \stage_1_retimer[7][14] , \stage_1_retimer[7][13] , 
        \stage_1_retimer[7][12] , \stage_1_retimer[7][11] , 
        \stage_1_retimer[7][10] , \stage_1_retimer[7][9] , 
        \stage_1_retimer[7][8] , \stage_1_retimer[7][7] , 
        \stage_1_retimer[7][6] , \stage_1_retimer[7][5] , 
        \stage_1_retimer[7][4] , \stage_1_retimer[7][3] , 
        \stage_1_retimer[7][2] , \stage_1_retimer[7][1] , 
        \stage_1_retimer[7][0] }), .in_control(in_control[8]), .out_upper({
        \stage_2_output[6][19] , \stage_2_output[6][18] , 
        \stage_2_output[6][17] , \stage_2_output[6][16] , 
        \stage_2_output[6][15] , \stage_2_output[6][14] , 
        \stage_2_output[6][13] , \stage_2_output[6][12] , 
        \stage_2_output[6][11] , \stage_2_output[6][10] , 
        \stage_2_output[6][9] , \stage_2_output[6][8] , \stage_2_output[6][7] , 
        \stage_2_output[6][6] , \stage_2_output[6][5] , \stage_2_output[6][4] , 
        \stage_2_output[6][3] , \stage_2_output[6][2] , \stage_2_output[6][1] , 
        \stage_2_output[6][0] }), .out_lower({\stage_2_output[7][19] , 
        \stage_2_output[7][18] , \stage_2_output[7][17] , 
        \stage_2_output[7][16] , \stage_2_output[7][15] , 
        \stage_2_output[7][14] , \stage_2_output[7][13] , 
        \stage_2_output[7][12] , \stage_2_output[7][11] , 
        \stage_2_output[7][10] , \stage_2_output[7][9] , 
        \stage_2_output[7][8] , \stage_2_output[7][7] , \stage_2_output[7][6] , 
        \stage_2_output[7][5] , \stage_2_output[7][4] , \stage_2_output[7][3] , 
        \stage_2_output[7][2] , \stage_2_output[7][1] , \stage_2_output[7][0] }) );
  crossbar_8 u_30_crossbar ( .in_upper({\stage_2_retimer[0][19] , 
        \stage_2_retimer[0][18] , \stage_2_retimer[0][17] , 
        \stage_2_retimer[0][16] , \stage_2_retimer[0][15] , 
        \stage_2_retimer[0][14] , \stage_2_retimer[0][13] , 
        \stage_2_retimer[0][12] , \stage_2_retimer[0][11] , 
        \stage_2_retimer[0][10] , \stage_2_retimer[0][9] , 
        \stage_2_retimer[0][8] , \stage_2_retimer[0][7] , 
        \stage_2_retimer[0][6] , \stage_2_retimer[0][5] , 
        \stage_2_retimer[0][4] , \stage_2_retimer[0][3] , 
        \stage_2_retimer[0][2] , \stage_2_retimer[0][1] , 
        \stage_2_retimer[0][0] }), .in_lower({\stage_2_retimer[2][19] , 
        \stage_2_retimer[2][18] , \stage_2_retimer[2][17] , 
        \stage_2_retimer[2][16] , \stage_2_retimer[2][15] , 
        \stage_2_retimer[2][14] , \stage_2_retimer[2][13] , 
        \stage_2_retimer[2][12] , \stage_2_retimer[2][11] , 
        \stage_2_retimer[2][10] , \stage_2_retimer[2][9] , 
        \stage_2_retimer[2][8] , \stage_2_retimer[2][7] , 
        \stage_2_retimer[2][6] , \stage_2_retimer[2][5] , 
        \stage_2_retimer[2][4] , \stage_2_retimer[2][3] , 
        \stage_2_retimer[2][2] , \stage_2_retimer[2][1] , 
        \stage_2_retimer[2][0] }), .in_control(in_control[7]), .out_upper({
        \stage_3_output[0][19] , \stage_3_output[0][18] , 
        \stage_3_output[0][17] , \stage_3_output[0][16] , 
        \stage_3_output[0][15] , \stage_3_output[0][14] , 
        \stage_3_output[0][13] , \stage_3_output[0][12] , 
        \stage_3_output[0][11] , \stage_3_output[0][10] , 
        \stage_3_output[0][9] , \stage_3_output[0][8] , \stage_3_output[0][7] , 
        \stage_3_output[0][6] , \stage_3_output[0][5] , \stage_3_output[0][4] , 
        \stage_3_output[0][3] , \stage_3_output[0][2] , \stage_3_output[0][1] , 
        \stage_3_output[0][0] }), .out_lower({\stage_3_output[1][19] , 
        \stage_3_output[1][18] , \stage_3_output[1][17] , 
        \stage_3_output[1][16] , \stage_3_output[1][15] , 
        \stage_3_output[1][14] , \stage_3_output[1][13] , 
        \stage_3_output[1][12] , \stage_3_output[1][11] , 
        \stage_3_output[1][10] , \stage_3_output[1][9] , 
        \stage_3_output[1][8] , \stage_3_output[1][7] , \stage_3_output[1][6] , 
        \stage_3_output[1][5] , \stage_3_output[1][4] , \stage_3_output[1][3] , 
        \stage_3_output[1][2] , \stage_3_output[1][1] , \stage_3_output[1][0] }) );
  crossbar_7 u_31_crossbar ( .in_upper({\stage_2_retimer[1][19] , 
        \stage_2_retimer[1][18] , \stage_2_retimer[1][17] , 
        \stage_2_retimer[1][16] , \stage_2_retimer[1][15] , 
        \stage_2_retimer[1][14] , \stage_2_retimer[1][13] , 
        \stage_2_retimer[1][12] , \stage_2_retimer[1][11] , 
        \stage_2_retimer[1][10] , \stage_2_retimer[1][9] , 
        \stage_2_retimer[1][8] , \stage_2_retimer[1][7] , 
        \stage_2_retimer[1][6] , \stage_2_retimer[1][5] , 
        \stage_2_retimer[1][4] , \stage_2_retimer[1][3] , 
        \stage_2_retimer[1][2] , \stage_2_retimer[1][1] , 
        \stage_2_retimer[1][0] }), .in_lower({\stage_2_retimer[3][19] , 
        \stage_2_retimer[3][18] , \stage_2_retimer[3][17] , 
        \stage_2_retimer[3][16] , \stage_2_retimer[3][15] , 
        \stage_2_retimer[3][14] , \stage_2_retimer[3][13] , 
        \stage_2_retimer[3][12] , \stage_2_retimer[3][11] , 
        \stage_2_retimer[3][10] , \stage_2_retimer[3][9] , 
        \stage_2_retimer[3][8] , \stage_2_retimer[3][7] , 
        \stage_2_retimer[3][6] , \stage_2_retimer[3][5] , 
        \stage_2_retimer[3][4] , \stage_2_retimer[3][3] , 
        \stage_2_retimer[3][2] , \stage_2_retimer[3][1] , 
        \stage_2_retimer[3][0] }), .in_control(in_control[6]), .out_upper({
        \stage_3_output[2][19] , \stage_3_output[2][18] , 
        \stage_3_output[2][17] , \stage_3_output[2][16] , 
        \stage_3_output[2][15] , \stage_3_output[2][14] , 
        \stage_3_output[2][13] , \stage_3_output[2][12] , 
        \stage_3_output[2][11] , \stage_3_output[2][10] , 
        \stage_3_output[2][9] , \stage_3_output[2][8] , \stage_3_output[2][7] , 
        \stage_3_output[2][6] , \stage_3_output[2][5] , \stage_3_output[2][4] , 
        \stage_3_output[2][3] , \stage_3_output[2][2] , \stage_3_output[2][1] , 
        \stage_3_output[2][0] }), .out_lower({\stage_3_output[3][19] , 
        \stage_3_output[3][18] , \stage_3_output[3][17] , 
        \stage_3_output[3][16] , \stage_3_output[3][15] , 
        \stage_3_output[3][14] , \stage_3_output[3][13] , 
        \stage_3_output[3][12] , \stage_3_output[3][11] , 
        \stage_3_output[3][10] , \stage_3_output[3][9] , 
        \stage_3_output[3][8] , \stage_3_output[3][7] , \stage_3_output[3][6] , 
        \stage_3_output[3][5] , \stage_3_output[3][4] , \stage_3_output[3][3] , 
        \stage_3_output[3][2] , \stage_3_output[3][1] , \stage_3_output[3][0] }) );
  crossbar_6 u_32_crossbar ( .in_upper({\stage_2_retimer[4][19] , 
        \stage_2_retimer[4][18] , \stage_2_retimer[4][17] , 
        \stage_2_retimer[4][16] , \stage_2_retimer[4][15] , 
        \stage_2_retimer[4][14] , \stage_2_retimer[4][13] , 
        \stage_2_retimer[4][12] , \stage_2_retimer[4][11] , 
        \stage_2_retimer[4][10] , \stage_2_retimer[4][9] , 
        \stage_2_retimer[4][8] , \stage_2_retimer[4][7] , 
        \stage_2_retimer[4][6] , \stage_2_retimer[4][5] , 
        \stage_2_retimer[4][4] , \stage_2_retimer[4][3] , 
        \stage_2_retimer[4][2] , \stage_2_retimer[4][1] , 
        \stage_2_retimer[4][0] }), .in_lower({\stage_2_retimer[6][19] , 
        \stage_2_retimer[6][18] , \stage_2_retimer[6][17] , 
        \stage_2_retimer[6][16] , \stage_2_retimer[6][15] , 
        \stage_2_retimer[6][14] , \stage_2_retimer[6][13] , 
        \stage_2_retimer[6][12] , \stage_2_retimer[6][11] , 
        \stage_2_retimer[6][10] , \stage_2_retimer[6][9] , 
        \stage_2_retimer[6][8] , \stage_2_retimer[6][7] , 
        \stage_2_retimer[6][6] , \stage_2_retimer[6][5] , 
        \stage_2_retimer[6][4] , \stage_2_retimer[6][3] , 
        \stage_2_retimer[6][2] , \stage_2_retimer[6][1] , 
        \stage_2_retimer[6][0] }), .in_control(in_control[5]), .out_upper({
        \stage_3_output[4][19] , \stage_3_output[4][18] , 
        \stage_3_output[4][17] , \stage_3_output[4][16] , 
        \stage_3_output[4][15] , \stage_3_output[4][14] , 
        \stage_3_output[4][13] , \stage_3_output[4][12] , 
        \stage_3_output[4][11] , \stage_3_output[4][10] , 
        \stage_3_output[4][9] , \stage_3_output[4][8] , \stage_3_output[4][7] , 
        \stage_3_output[4][6] , \stage_3_output[4][5] , \stage_3_output[4][4] , 
        \stage_3_output[4][3] , \stage_3_output[4][2] , \stage_3_output[4][1] , 
        \stage_3_output[4][0] }), .out_lower({\stage_3_output[5][19] , 
        \stage_3_output[5][18] , \stage_3_output[5][17] , 
        \stage_3_output[5][16] , \stage_3_output[5][15] , 
        \stage_3_output[5][14] , \stage_3_output[5][13] , 
        \stage_3_output[5][12] , \stage_3_output[5][11] , 
        \stage_3_output[5][10] , \stage_3_output[5][9] , 
        \stage_3_output[5][8] , \stage_3_output[5][7] , \stage_3_output[5][6] , 
        \stage_3_output[5][5] , \stage_3_output[5][4] , \stage_3_output[5][3] , 
        \stage_3_output[5][2] , \stage_3_output[5][1] , \stage_3_output[5][0] }) );
  crossbar_5 u_33_crossbar ( .in_upper({\stage_2_retimer[5][19] , 
        \stage_2_retimer[5][18] , \stage_2_retimer[5][17] , 
        \stage_2_retimer[5][16] , \stage_2_retimer[5][15] , 
        \stage_2_retimer[5][14] , \stage_2_retimer[5][13] , 
        \stage_2_retimer[5][12] , \stage_2_retimer[5][11] , 
        \stage_2_retimer[5][10] , \stage_2_retimer[5][9] , 
        \stage_2_retimer[5][8] , \stage_2_retimer[5][7] , 
        \stage_2_retimer[5][6] , \stage_2_retimer[5][5] , 
        \stage_2_retimer[5][4] , \stage_2_retimer[5][3] , 
        \stage_2_retimer[5][2] , \stage_2_retimer[5][1] , 
        \stage_2_retimer[5][0] }), .in_lower({\stage_2_retimer[7][19] , 
        \stage_2_retimer[7][18] , \stage_2_retimer[7][17] , 
        \stage_2_retimer[7][16] , \stage_2_retimer[7][15] , 
        \stage_2_retimer[7][14] , \stage_2_retimer[7][13] , 
        \stage_2_retimer[7][12] , \stage_2_retimer[7][11] , 
        \stage_2_retimer[7][10] , \stage_2_retimer[7][9] , 
        \stage_2_retimer[7][8] , \stage_2_retimer[7][7] , 
        \stage_2_retimer[7][6] , \stage_2_retimer[7][5] , 
        \stage_2_retimer[7][4] , \stage_2_retimer[7][3] , 
        \stage_2_retimer[7][2] , \stage_2_retimer[7][1] , 
        \stage_2_retimer[7][0] }), .in_control(in_control[4]), .out_upper({
        \stage_3_output[6][19] , \stage_3_output[6][18] , 
        \stage_3_output[6][17] , \stage_3_output[6][16] , 
        \stage_3_output[6][15] , \stage_3_output[6][14] , 
        \stage_3_output[6][13] , \stage_3_output[6][12] , 
        \stage_3_output[6][11] , \stage_3_output[6][10] , 
        \stage_3_output[6][9] , \stage_3_output[6][8] , \stage_3_output[6][7] , 
        \stage_3_output[6][6] , \stage_3_output[6][5] , \stage_3_output[6][4] , 
        \stage_3_output[6][3] , \stage_3_output[6][2] , \stage_3_output[6][1] , 
        \stage_3_output[6][0] }), .out_lower({\stage_3_output[7][19] , 
        \stage_3_output[7][18] , \stage_3_output[7][17] , 
        \stage_3_output[7][16] , \stage_3_output[7][15] , 
        \stage_3_output[7][14] , \stage_3_output[7][13] , 
        \stage_3_output[7][12] , \stage_3_output[7][11] , 
        \stage_3_output[7][10] , \stage_3_output[7][9] , 
        \stage_3_output[7][8] , \stage_3_output[7][7] , \stage_3_output[7][6] , 
        \stage_3_output[7][5] , \stage_3_output[7][4] , \stage_3_output[7][3] , 
        \stage_3_output[7][2] , \stage_3_output[7][1] , \stage_3_output[7][0] }) );
  crossbar_4 u_40_crossbar ( .in_upper({\stage_3_retimer[0][19] , 
        \stage_3_retimer[0][18] , \stage_3_retimer[0][17] , 
        \stage_3_retimer[0][16] , \stage_3_retimer[0][15] , 
        \stage_3_retimer[0][14] , \stage_3_retimer[0][13] , 
        \stage_3_retimer[0][12] , \stage_3_retimer[0][11] , 
        \stage_3_retimer[0][10] , \stage_3_retimer[0][9] , 
        \stage_3_retimer[0][8] , \stage_3_retimer[0][7] , 
        \stage_3_retimer[0][6] , \stage_3_retimer[0][5] , 
        \stage_3_retimer[0][4] , \stage_3_retimer[0][3] , 
        \stage_3_retimer[0][2] , \stage_3_retimer[0][1] , 
        \stage_3_retimer[0][0] }), .in_lower({\stage_3_retimer[4][19] , 
        \stage_3_retimer[4][18] , \stage_3_retimer[4][17] , 
        \stage_3_retimer[4][16] , \stage_3_retimer[4][15] , 
        \stage_3_retimer[4][14] , \stage_3_retimer[4][13] , 
        \stage_3_retimer[4][12] , \stage_3_retimer[4][11] , 
        \stage_3_retimer[4][10] , \stage_3_retimer[4][9] , 
        \stage_3_retimer[4][8] , \stage_3_retimer[4][7] , 
        \stage_3_retimer[4][6] , \stage_3_retimer[4][5] , 
        \stage_3_retimer[4][4] , \stage_3_retimer[4][3] , 
        \stage_3_retimer[4][2] , \stage_3_retimer[4][1] , 
        \stage_3_retimer[4][0] }), .in_control(in_control[3]), .out_upper({
        \stage_4_output[0][19] , \stage_4_output[0][18] , 
        \stage_4_output[0][17] , \stage_4_output[0][16] , 
        \stage_4_output[0][15] , \stage_4_output[0][14] , 
        \stage_4_output[0][13] , \stage_4_output[0][12] , 
        \stage_4_output[0][11] , \stage_4_output[0][10] , 
        \stage_4_output[0][9] , \stage_4_output[0][8] , \stage_4_output[0][7] , 
        \stage_4_output[0][6] , \stage_4_output[0][5] , \stage_4_output[0][4] , 
        \stage_4_output[0][3] , \stage_4_output[0][2] , \stage_4_output[0][1] , 
        \stage_4_output[0][0] }), .out_lower({\stage_4_output[1][19] , 
        \stage_4_output[1][18] , \stage_4_output[1][17] , 
        \stage_4_output[1][16] , \stage_4_output[1][15] , 
        \stage_4_output[1][14] , \stage_4_output[1][13] , 
        \stage_4_output[1][12] , \stage_4_output[1][11] , 
        \stage_4_output[1][10] , \stage_4_output[1][9] , 
        \stage_4_output[1][8] , \stage_4_output[1][7] , \stage_4_output[1][6] , 
        \stage_4_output[1][5] , \stage_4_output[1][4] , \stage_4_output[1][3] , 
        \stage_4_output[1][2] , \stage_4_output[1][1] , \stage_4_output[1][0] }) );
  crossbar_3 u_41_crossbar ( .in_upper({\stage_3_retimer[1][19] , 
        \stage_3_retimer[1][18] , \stage_3_retimer[1][17] , 
        \stage_3_retimer[1][16] , \stage_3_retimer[1][15] , 
        \stage_3_retimer[1][14] , \stage_3_retimer[1][13] , 
        \stage_3_retimer[1][12] , \stage_3_retimer[1][11] , 
        \stage_3_retimer[1][10] , \stage_3_retimer[1][9] , 
        \stage_3_retimer[1][8] , \stage_3_retimer[1][7] , 
        \stage_3_retimer[1][6] , \stage_3_retimer[1][5] , 
        \stage_3_retimer[1][4] , \stage_3_retimer[1][3] , 
        \stage_3_retimer[1][2] , \stage_3_retimer[1][1] , 
        \stage_3_retimer[1][0] }), .in_lower({\stage_3_retimer[5][19] , 
        \stage_3_retimer[5][18] , \stage_3_retimer[5][17] , 
        \stage_3_retimer[5][16] , \stage_3_retimer[5][15] , 
        \stage_3_retimer[5][14] , \stage_3_retimer[5][13] , 
        \stage_3_retimer[5][12] , \stage_3_retimer[5][11] , 
        \stage_3_retimer[5][10] , \stage_3_retimer[5][9] , 
        \stage_3_retimer[5][8] , \stage_3_retimer[5][7] , 
        \stage_3_retimer[5][6] , \stage_3_retimer[5][5] , 
        \stage_3_retimer[5][4] , \stage_3_retimer[5][3] , 
        \stage_3_retimer[5][2] , \stage_3_retimer[5][1] , 
        \stage_3_retimer[5][0] }), .in_control(in_control[2]), .out_upper({
        \stage_4_output[2][19] , \stage_4_output[2][18] , 
        \stage_4_output[2][17] , \stage_4_output[2][16] , 
        \stage_4_output[2][15] , \stage_4_output[2][14] , 
        \stage_4_output[2][13] , \stage_4_output[2][12] , 
        \stage_4_output[2][11] , \stage_4_output[2][10] , 
        \stage_4_output[2][9] , \stage_4_output[2][8] , \stage_4_output[2][7] , 
        \stage_4_output[2][6] , \stage_4_output[2][5] , \stage_4_output[2][4] , 
        \stage_4_output[2][3] , \stage_4_output[2][2] , \stage_4_output[2][1] , 
        \stage_4_output[2][0] }), .out_lower({\stage_4_output[3][19] , 
        \stage_4_output[3][18] , \stage_4_output[3][17] , 
        \stage_4_output[3][16] , \stage_4_output[3][15] , 
        \stage_4_output[3][14] , \stage_4_output[3][13] , 
        \stage_4_output[3][12] , \stage_4_output[3][11] , 
        \stage_4_output[3][10] , \stage_4_output[3][9] , 
        \stage_4_output[3][8] , \stage_4_output[3][7] , \stage_4_output[3][6] , 
        \stage_4_output[3][5] , \stage_4_output[3][4] , \stage_4_output[3][3] , 
        \stage_4_output[3][2] , \stage_4_output[3][1] , \stage_4_output[3][0] }) );
  crossbar_2 u_42_crossbar ( .in_upper({\stage_3_retimer[2][19] , 
        \stage_3_retimer[2][18] , \stage_3_retimer[2][17] , 
        \stage_3_retimer[2][16] , \stage_3_retimer[2][15] , 
        \stage_3_retimer[2][14] , \stage_3_retimer[2][13] , 
        \stage_3_retimer[2][12] , \stage_3_retimer[2][11] , 
        \stage_3_retimer[2][10] , \stage_3_retimer[2][9] , 
        \stage_3_retimer[2][8] , \stage_3_retimer[2][7] , 
        \stage_3_retimer[2][6] , \stage_3_retimer[2][5] , 
        \stage_3_retimer[2][4] , \stage_3_retimer[2][3] , 
        \stage_3_retimer[2][2] , \stage_3_retimer[2][1] , 
        \stage_3_retimer[2][0] }), .in_lower({\stage_3_retimer[6][19] , 
        \stage_3_retimer[6][18] , \stage_3_retimer[6][17] , 
        \stage_3_retimer[6][16] , \stage_3_retimer[6][15] , 
        \stage_3_retimer[6][14] , \stage_3_retimer[6][13] , 
        \stage_3_retimer[6][12] , \stage_3_retimer[6][11] , 
        \stage_3_retimer[6][10] , \stage_3_retimer[6][9] , 
        \stage_3_retimer[6][8] , \stage_3_retimer[6][7] , 
        \stage_3_retimer[6][6] , \stage_3_retimer[6][5] , 
        \stage_3_retimer[6][4] , \stage_3_retimer[6][3] , 
        \stage_3_retimer[6][2] , \stage_3_retimer[6][1] , 
        \stage_3_retimer[6][0] }), .in_control(in_control[1]), .out_upper({
        \stage_4_output[4][19] , \stage_4_output[4][18] , 
        \stage_4_output[4][17] , \stage_4_output[4][16] , 
        \stage_4_output[4][15] , \stage_4_output[4][14] , 
        \stage_4_output[4][13] , \stage_4_output[4][12] , 
        \stage_4_output[4][11] , \stage_4_output[4][10] , 
        \stage_4_output[4][9] , \stage_4_output[4][8] , \stage_4_output[4][7] , 
        \stage_4_output[4][6] , \stage_4_output[4][5] , \stage_4_output[4][4] , 
        \stage_4_output[4][3] , \stage_4_output[4][2] , \stage_4_output[4][1] , 
        \stage_4_output[4][0] }), .out_lower({\stage_4_output[5][19] , 
        \stage_4_output[5][18] , \stage_4_output[5][17] , 
        \stage_4_output[5][16] , \stage_4_output[5][15] , 
        \stage_4_output[5][14] , \stage_4_output[5][13] , 
        \stage_4_output[5][12] , \stage_4_output[5][11] , 
        \stage_4_output[5][10] , \stage_4_output[5][9] , 
        \stage_4_output[5][8] , \stage_4_output[5][7] , \stage_4_output[5][6] , 
        \stage_4_output[5][5] , \stage_4_output[5][4] , \stage_4_output[5][3] , 
        \stage_4_output[5][2] , \stage_4_output[5][1] , \stage_4_output[5][0] }) );
  crossbar_1 u_43_crossbar ( .in_upper({\stage_3_retimer[3][19] , 
        \stage_3_retimer[3][18] , \stage_3_retimer[3][17] , 
        \stage_3_retimer[3][16] , \stage_3_retimer[3][15] , 
        \stage_3_retimer[3][14] , \stage_3_retimer[3][13] , 
        \stage_3_retimer[3][12] , \stage_3_retimer[3][11] , 
        \stage_3_retimer[3][10] , \stage_3_retimer[3][9] , 
        \stage_3_retimer[3][8] , \stage_3_retimer[3][7] , 
        \stage_3_retimer[3][6] , \stage_3_retimer[3][5] , 
        \stage_3_retimer[3][4] , \stage_3_retimer[3][3] , 
        \stage_3_retimer[3][2] , \stage_3_retimer[3][1] , 
        \stage_3_retimer[3][0] }), .in_lower({\stage_3_retimer[7][19] , 
        \stage_3_retimer[7][18] , \stage_3_retimer[7][17] , 
        \stage_3_retimer[7][16] , \stage_3_retimer[7][15] , 
        \stage_3_retimer[7][14] , \stage_3_retimer[7][13] , 
        \stage_3_retimer[7][12] , \stage_3_retimer[7][11] , 
        \stage_3_retimer[7][10] , \stage_3_retimer[7][9] , 
        \stage_3_retimer[7][8] , \stage_3_retimer[7][7] , 
        \stage_3_retimer[7][6] , \stage_3_retimer[7][5] , 
        \stage_3_retimer[7][4] , \stage_3_retimer[7][3] , 
        \stage_3_retimer[7][2] , \stage_3_retimer[7][1] , 
        \stage_3_retimer[7][0] }), .in_control(in_control[0]), .out_upper({
        \stage_4_output[6][19] , \stage_4_output[6][18] , 
        \stage_4_output[6][17] , \stage_4_output[6][16] , 
        \stage_4_output[6][15] , \stage_4_output[6][14] , 
        \stage_4_output[6][13] , \stage_4_output[6][12] , 
        \stage_4_output[6][11] , \stage_4_output[6][10] , 
        \stage_4_output[6][9] , \stage_4_output[6][8] , \stage_4_output[6][7] , 
        \stage_4_output[6][6] , \stage_4_output[6][5] , \stage_4_output[6][4] , 
        \stage_4_output[6][3] , \stage_4_output[6][2] , \stage_4_output[6][1] , 
        \stage_4_output[6][0] }), .out_lower({\stage_4_output[7][19] , 
        \stage_4_output[7][18] , \stage_4_output[7][17] , 
        \stage_4_output[7][16] , \stage_4_output[7][15] , 
        \stage_4_output[7][14] , \stage_4_output[7][13] , 
        \stage_4_output[7][12] , \stage_4_output[7][11] , 
        \stage_4_output[7][10] , \stage_4_output[7][9] , 
        \stage_4_output[7][8] , \stage_4_output[7][7] , \stage_4_output[7][6] , 
        \stage_4_output[7][5] , \stage_4_output[7][4] , \stage_4_output[7][3] , 
        \stage_4_output[7][2] , \stage_4_output[7][1] , \stage_4_output[7][0] }) );
  DFQD1 \stage_0_retimer_reg[7][19]  ( .D(\stage_0_output[7][19] ), .CP(clk), 
        .Q(\stage_0_retimer[7][19] ) );
  DFQD1 \stage_0_retimer_reg[7][18]  ( .D(\stage_0_output[7][18] ), .CP(clk), 
        .Q(\stage_0_retimer[7][18] ) );
  DFQD1 \stage_0_retimer_reg[7][17]  ( .D(\stage_0_output[7][17] ), .CP(clk), 
        .Q(\stage_0_retimer[7][17] ) );
  DFQD1 \stage_0_retimer_reg[7][16]  ( .D(\stage_0_output[7][16] ), .CP(clk), 
        .Q(\stage_0_retimer[7][16] ) );
  DFQD1 \stage_0_retimer_reg[7][15]  ( .D(\stage_0_output[7][15] ), .CP(clk), 
        .Q(\stage_0_retimer[7][15] ) );
  DFQD1 \stage_0_retimer_reg[7][14]  ( .D(\stage_0_output[7][14] ), .CP(clk), 
        .Q(\stage_0_retimer[7][14] ) );
  DFQD1 \stage_0_retimer_reg[7][13]  ( .D(\stage_0_output[7][13] ), .CP(clk), 
        .Q(\stage_0_retimer[7][13] ) );
  DFQD1 \stage_0_retimer_reg[7][12]  ( .D(\stage_0_output[7][12] ), .CP(clk), 
        .Q(\stage_0_retimer[7][12] ) );
  DFQD1 \stage_0_retimer_reg[7][11]  ( .D(\stage_0_output[7][11] ), .CP(clk), 
        .Q(\stage_0_retimer[7][11] ) );
  DFQD1 \stage_0_retimer_reg[7][10]  ( .D(\stage_0_output[7][10] ), .CP(clk), 
        .Q(\stage_0_retimer[7][10] ) );
  DFQD1 \stage_0_retimer_reg[7][9]  ( .D(\stage_0_output[7][9] ), .CP(clk), 
        .Q(\stage_0_retimer[7][9] ) );
  DFQD1 \stage_0_retimer_reg[7][8]  ( .D(\stage_0_output[7][8] ), .CP(clk), 
        .Q(\stage_0_retimer[7][8] ) );
  DFQD1 \stage_0_retimer_reg[7][7]  ( .D(\stage_0_output[7][7] ), .CP(clk), 
        .Q(\stage_0_retimer[7][7] ) );
  DFQD1 \stage_0_retimer_reg[7][6]  ( .D(\stage_0_output[7][6] ), .CP(clk), 
        .Q(\stage_0_retimer[7][6] ) );
  DFQD1 \stage_0_retimer_reg[7][5]  ( .D(\stage_0_output[7][5] ), .CP(clk), 
        .Q(\stage_0_retimer[7][5] ) );
  DFQD1 \stage_0_retimer_reg[7][4]  ( .D(\stage_0_output[7][4] ), .CP(clk), 
        .Q(\stage_0_retimer[7][4] ) );
  DFQD1 \stage_0_retimer_reg[7][3]  ( .D(\stage_0_output[7][3] ), .CP(clk), 
        .Q(\stage_0_retimer[7][3] ) );
  DFQD1 \stage_0_retimer_reg[7][2]  ( .D(\stage_0_output[7][2] ), .CP(clk), 
        .Q(\stage_0_retimer[7][2] ) );
  DFQD1 \stage_0_retimer_reg[7][1]  ( .D(\stage_0_output[7][1] ), .CP(clk), 
        .Q(\stage_0_retimer[7][1] ) );
  DFQD1 \stage_0_retimer_reg[7][0]  ( .D(\stage_0_output[7][0] ), .CP(clk), 
        .Q(\stage_0_retimer[7][0] ) );
  DFQD1 \stage_0_retimer_reg[6][19]  ( .D(\stage_0_output[6][19] ), .CP(clk), 
        .Q(\stage_0_retimer[6][19] ) );
  DFQD1 \stage_0_retimer_reg[6][18]  ( .D(\stage_0_output[6][18] ), .CP(clk), 
        .Q(\stage_0_retimer[6][18] ) );
  DFQD1 \stage_0_retimer_reg[6][17]  ( .D(\stage_0_output[6][17] ), .CP(clk), 
        .Q(\stage_0_retimer[6][17] ) );
  DFQD1 \stage_0_retimer_reg[6][16]  ( .D(\stage_0_output[6][16] ), .CP(clk), 
        .Q(\stage_0_retimer[6][16] ) );
  DFQD1 \stage_0_retimer_reg[6][15]  ( .D(\stage_0_output[6][15] ), .CP(clk), 
        .Q(\stage_0_retimer[6][15] ) );
  DFQD1 \stage_0_retimer_reg[6][14]  ( .D(\stage_0_output[6][14] ), .CP(clk), 
        .Q(\stage_0_retimer[6][14] ) );
  DFQD1 \stage_0_retimer_reg[6][13]  ( .D(\stage_0_output[6][13] ), .CP(clk), 
        .Q(\stage_0_retimer[6][13] ) );
  DFQD1 \stage_0_retimer_reg[6][12]  ( .D(\stage_0_output[6][12] ), .CP(clk), 
        .Q(\stage_0_retimer[6][12] ) );
  DFQD1 \stage_0_retimer_reg[6][11]  ( .D(\stage_0_output[6][11] ), .CP(clk), 
        .Q(\stage_0_retimer[6][11] ) );
  DFQD1 \stage_0_retimer_reg[6][10]  ( .D(\stage_0_output[6][10] ), .CP(clk), 
        .Q(\stage_0_retimer[6][10] ) );
  DFQD1 \stage_0_retimer_reg[6][9]  ( .D(\stage_0_output[6][9] ), .CP(clk), 
        .Q(\stage_0_retimer[6][9] ) );
  DFQD1 \stage_0_retimer_reg[6][8]  ( .D(\stage_0_output[6][8] ), .CP(clk), 
        .Q(\stage_0_retimer[6][8] ) );
  DFQD1 \stage_0_retimer_reg[6][7]  ( .D(\stage_0_output[6][7] ), .CP(clk), 
        .Q(\stage_0_retimer[6][7] ) );
  DFQD1 \stage_0_retimer_reg[6][6]  ( .D(\stage_0_output[6][6] ), .CP(clk), 
        .Q(\stage_0_retimer[6][6] ) );
  DFQD1 \stage_0_retimer_reg[6][5]  ( .D(\stage_0_output[6][5] ), .CP(clk), 
        .Q(\stage_0_retimer[6][5] ) );
  DFQD1 \stage_0_retimer_reg[6][4]  ( .D(\stage_0_output[6][4] ), .CP(clk), 
        .Q(\stage_0_retimer[6][4] ) );
  DFQD1 \stage_0_retimer_reg[6][3]  ( .D(\stage_0_output[6][3] ), .CP(clk), 
        .Q(\stage_0_retimer[6][3] ) );
  DFQD1 \stage_0_retimer_reg[6][2]  ( .D(\stage_0_output[6][2] ), .CP(clk), 
        .Q(\stage_0_retimer[6][2] ) );
  DFQD1 \stage_0_retimer_reg[6][1]  ( .D(\stage_0_output[6][1] ), .CP(clk), 
        .Q(\stage_0_retimer[6][1] ) );
  DFQD1 \stage_0_retimer_reg[6][0]  ( .D(\stage_0_output[6][0] ), .CP(clk), 
        .Q(\stage_0_retimer[6][0] ) );
  DFQD1 \stage_0_retimer_reg[5][19]  ( .D(\stage_0_output[5][19] ), .CP(clk), 
        .Q(\stage_0_retimer[5][19] ) );
  DFQD1 \stage_0_retimer_reg[5][18]  ( .D(\stage_0_output[5][18] ), .CP(clk), 
        .Q(\stage_0_retimer[5][18] ) );
  DFQD1 \stage_0_retimer_reg[5][17]  ( .D(\stage_0_output[5][17] ), .CP(clk), 
        .Q(\stage_0_retimer[5][17] ) );
  DFQD1 \stage_0_retimer_reg[5][16]  ( .D(\stage_0_output[5][16] ), .CP(clk), 
        .Q(\stage_0_retimer[5][16] ) );
  DFQD1 \stage_0_retimer_reg[5][15]  ( .D(\stage_0_output[5][15] ), .CP(clk), 
        .Q(\stage_0_retimer[5][15] ) );
  DFQD1 \stage_0_retimer_reg[5][14]  ( .D(\stage_0_output[5][14] ), .CP(clk), 
        .Q(\stage_0_retimer[5][14] ) );
  DFQD1 \stage_0_retimer_reg[5][13]  ( .D(\stage_0_output[5][13] ), .CP(clk), 
        .Q(\stage_0_retimer[5][13] ) );
  DFQD1 \stage_0_retimer_reg[5][12]  ( .D(\stage_0_output[5][12] ), .CP(clk), 
        .Q(\stage_0_retimer[5][12] ) );
  DFQD1 \stage_0_retimer_reg[5][11]  ( .D(\stage_0_output[5][11] ), .CP(clk), 
        .Q(\stage_0_retimer[5][11] ) );
  DFQD1 \stage_0_retimer_reg[5][10]  ( .D(\stage_0_output[5][10] ), .CP(clk), 
        .Q(\stage_0_retimer[5][10] ) );
  DFQD1 \stage_0_retimer_reg[5][9]  ( .D(\stage_0_output[5][9] ), .CP(clk), 
        .Q(\stage_0_retimer[5][9] ) );
  DFQD1 \stage_0_retimer_reg[5][8]  ( .D(\stage_0_output[5][8] ), .CP(clk), 
        .Q(\stage_0_retimer[5][8] ) );
  DFQD1 \stage_0_retimer_reg[5][7]  ( .D(\stage_0_output[5][7] ), .CP(clk), 
        .Q(\stage_0_retimer[5][7] ) );
  DFQD1 \stage_0_retimer_reg[5][6]  ( .D(\stage_0_output[5][6] ), .CP(clk), 
        .Q(\stage_0_retimer[5][6] ) );
  DFQD1 \stage_0_retimer_reg[5][5]  ( .D(\stage_0_output[5][5] ), .CP(clk), 
        .Q(\stage_0_retimer[5][5] ) );
  DFQD1 \stage_0_retimer_reg[5][4]  ( .D(\stage_0_output[5][4] ), .CP(clk), 
        .Q(\stage_0_retimer[5][4] ) );
  DFQD1 \stage_0_retimer_reg[5][3]  ( .D(\stage_0_output[5][3] ), .CP(clk), 
        .Q(\stage_0_retimer[5][3] ) );
  DFQD1 \stage_0_retimer_reg[5][2]  ( .D(\stage_0_output[5][2] ), .CP(clk), 
        .Q(\stage_0_retimer[5][2] ) );
  DFQD1 \stage_0_retimer_reg[5][1]  ( .D(\stage_0_output[5][1] ), .CP(clk), 
        .Q(\stage_0_retimer[5][1] ) );
  DFQD1 \stage_0_retimer_reg[5][0]  ( .D(\stage_0_output[5][0] ), .CP(clk), 
        .Q(\stage_0_retimer[5][0] ) );
  DFQD1 \stage_0_retimer_reg[4][19]  ( .D(\stage_0_output[4][19] ), .CP(clk), 
        .Q(\stage_0_retimer[4][19] ) );
  DFQD1 \stage_0_retimer_reg[4][18]  ( .D(\stage_0_output[4][18] ), .CP(clk), 
        .Q(\stage_0_retimer[4][18] ) );
  DFQD1 \stage_0_retimer_reg[4][17]  ( .D(\stage_0_output[4][17] ), .CP(clk), 
        .Q(\stage_0_retimer[4][17] ) );
  DFQD1 \stage_0_retimer_reg[4][16]  ( .D(\stage_0_output[4][16] ), .CP(clk), 
        .Q(\stage_0_retimer[4][16] ) );
  DFQD1 \stage_0_retimer_reg[4][15]  ( .D(\stage_0_output[4][15] ), .CP(clk), 
        .Q(\stage_0_retimer[4][15] ) );
  DFQD1 \stage_0_retimer_reg[4][14]  ( .D(\stage_0_output[4][14] ), .CP(clk), 
        .Q(\stage_0_retimer[4][14] ) );
  DFQD1 \stage_0_retimer_reg[4][13]  ( .D(\stage_0_output[4][13] ), .CP(clk), 
        .Q(\stage_0_retimer[4][13] ) );
  DFQD1 \stage_0_retimer_reg[4][12]  ( .D(\stage_0_output[4][12] ), .CP(clk), 
        .Q(\stage_0_retimer[4][12] ) );
  DFQD1 \stage_0_retimer_reg[4][11]  ( .D(\stage_0_output[4][11] ), .CP(clk), 
        .Q(\stage_0_retimer[4][11] ) );
  DFQD1 \stage_0_retimer_reg[4][10]  ( .D(\stage_0_output[4][10] ), .CP(clk), 
        .Q(\stage_0_retimer[4][10] ) );
  DFQD1 \stage_0_retimer_reg[4][9]  ( .D(\stage_0_output[4][9] ), .CP(clk), 
        .Q(\stage_0_retimer[4][9] ) );
  DFQD1 \stage_0_retimer_reg[4][8]  ( .D(\stage_0_output[4][8] ), .CP(clk), 
        .Q(\stage_0_retimer[4][8] ) );
  DFQD1 \stage_0_retimer_reg[4][7]  ( .D(\stage_0_output[4][7] ), .CP(clk), 
        .Q(\stage_0_retimer[4][7] ) );
  DFQD1 \stage_0_retimer_reg[4][6]  ( .D(\stage_0_output[4][6] ), .CP(clk), 
        .Q(\stage_0_retimer[4][6] ) );
  DFQD1 \stage_0_retimer_reg[4][5]  ( .D(\stage_0_output[4][5] ), .CP(clk), 
        .Q(\stage_0_retimer[4][5] ) );
  DFQD1 \stage_0_retimer_reg[4][4]  ( .D(\stage_0_output[4][4] ), .CP(clk), 
        .Q(\stage_0_retimer[4][4] ) );
  DFQD1 \stage_0_retimer_reg[4][3]  ( .D(\stage_0_output[4][3] ), .CP(clk), 
        .Q(\stage_0_retimer[4][3] ) );
  DFQD1 \stage_0_retimer_reg[4][2]  ( .D(\stage_0_output[4][2] ), .CP(clk), 
        .Q(\stage_0_retimer[4][2] ) );
  DFQD1 \stage_0_retimer_reg[4][1]  ( .D(\stage_0_output[4][1] ), .CP(clk), 
        .Q(\stage_0_retimer[4][1] ) );
  DFQD1 \stage_0_retimer_reg[4][0]  ( .D(\stage_0_output[4][0] ), .CP(clk), 
        .Q(\stage_0_retimer[4][0] ) );
  DFQD1 \stage_0_retimer_reg[3][19]  ( .D(\stage_0_output[3][19] ), .CP(clk), 
        .Q(\stage_0_retimer[3][19] ) );
  DFQD1 \stage_0_retimer_reg[3][18]  ( .D(\stage_0_output[3][18] ), .CP(clk), 
        .Q(\stage_0_retimer[3][18] ) );
  DFQD1 \stage_0_retimer_reg[3][17]  ( .D(\stage_0_output[3][17] ), .CP(clk), 
        .Q(\stage_0_retimer[3][17] ) );
  DFQD1 \stage_0_retimer_reg[3][16]  ( .D(\stage_0_output[3][16] ), .CP(clk), 
        .Q(\stage_0_retimer[3][16] ) );
  DFQD1 \stage_0_retimer_reg[3][15]  ( .D(\stage_0_output[3][15] ), .CP(clk), 
        .Q(\stage_0_retimer[3][15] ) );
  DFQD1 \stage_0_retimer_reg[3][14]  ( .D(\stage_0_output[3][14] ), .CP(clk), 
        .Q(\stage_0_retimer[3][14] ) );
  DFQD1 \stage_0_retimer_reg[3][13]  ( .D(\stage_0_output[3][13] ), .CP(clk), 
        .Q(\stage_0_retimer[3][13] ) );
  DFQD1 \stage_0_retimer_reg[3][12]  ( .D(\stage_0_output[3][12] ), .CP(clk), 
        .Q(\stage_0_retimer[3][12] ) );
  DFQD1 \stage_0_retimer_reg[3][11]  ( .D(\stage_0_output[3][11] ), .CP(clk), 
        .Q(\stage_0_retimer[3][11] ) );
  DFQD1 \stage_0_retimer_reg[3][10]  ( .D(\stage_0_output[3][10] ), .CP(clk), 
        .Q(\stage_0_retimer[3][10] ) );
  DFQD1 \stage_0_retimer_reg[3][9]  ( .D(\stage_0_output[3][9] ), .CP(clk), 
        .Q(\stage_0_retimer[3][9] ) );
  DFQD1 \stage_0_retimer_reg[3][8]  ( .D(\stage_0_output[3][8] ), .CP(clk), 
        .Q(\stage_0_retimer[3][8] ) );
  DFQD1 \stage_0_retimer_reg[3][7]  ( .D(\stage_0_output[3][7] ), .CP(clk), 
        .Q(\stage_0_retimer[3][7] ) );
  DFQD1 \stage_0_retimer_reg[3][6]  ( .D(\stage_0_output[3][6] ), .CP(clk), 
        .Q(\stage_0_retimer[3][6] ) );
  DFQD1 \stage_0_retimer_reg[3][5]  ( .D(\stage_0_output[3][5] ), .CP(clk), 
        .Q(\stage_0_retimer[3][5] ) );
  DFQD1 \stage_0_retimer_reg[3][4]  ( .D(\stage_0_output[3][4] ), .CP(clk), 
        .Q(\stage_0_retimer[3][4] ) );
  DFQD1 \stage_0_retimer_reg[3][3]  ( .D(\stage_0_output[3][3] ), .CP(clk), 
        .Q(\stage_0_retimer[3][3] ) );
  DFQD1 \stage_0_retimer_reg[3][2]  ( .D(\stage_0_output[3][2] ), .CP(clk), 
        .Q(\stage_0_retimer[3][2] ) );
  DFQD1 \stage_0_retimer_reg[3][1]  ( .D(\stage_0_output[3][1] ), .CP(clk), 
        .Q(\stage_0_retimer[3][1] ) );
  DFQD1 \stage_0_retimer_reg[3][0]  ( .D(\stage_0_output[3][0] ), .CP(clk), 
        .Q(\stage_0_retimer[3][0] ) );
  DFQD1 \stage_0_retimer_reg[2][19]  ( .D(\stage_0_output[2][19] ), .CP(clk), 
        .Q(\stage_0_retimer[2][19] ) );
  DFQD1 \stage_0_retimer_reg[2][18]  ( .D(\stage_0_output[2][18] ), .CP(clk), 
        .Q(\stage_0_retimer[2][18] ) );
  DFQD1 \stage_0_retimer_reg[2][17]  ( .D(\stage_0_output[2][17] ), .CP(clk), 
        .Q(\stage_0_retimer[2][17] ) );
  DFQD1 \stage_0_retimer_reg[2][16]  ( .D(\stage_0_output[2][16] ), .CP(clk), 
        .Q(\stage_0_retimer[2][16] ) );
  DFQD1 \stage_0_retimer_reg[2][15]  ( .D(\stage_0_output[2][15] ), .CP(clk), 
        .Q(\stage_0_retimer[2][15] ) );
  DFQD1 \stage_0_retimer_reg[2][14]  ( .D(\stage_0_output[2][14] ), .CP(clk), 
        .Q(\stage_0_retimer[2][14] ) );
  DFQD1 \stage_0_retimer_reg[2][13]  ( .D(\stage_0_output[2][13] ), .CP(clk), 
        .Q(\stage_0_retimer[2][13] ) );
  DFQD1 \stage_0_retimer_reg[2][12]  ( .D(\stage_0_output[2][12] ), .CP(clk), 
        .Q(\stage_0_retimer[2][12] ) );
  DFQD1 \stage_0_retimer_reg[2][11]  ( .D(\stage_0_output[2][11] ), .CP(clk), 
        .Q(\stage_0_retimer[2][11] ) );
  DFQD1 \stage_0_retimer_reg[2][10]  ( .D(\stage_0_output[2][10] ), .CP(clk), 
        .Q(\stage_0_retimer[2][10] ) );
  DFQD1 \stage_0_retimer_reg[2][9]  ( .D(\stage_0_output[2][9] ), .CP(clk), 
        .Q(\stage_0_retimer[2][9] ) );
  DFQD1 \stage_0_retimer_reg[2][8]  ( .D(\stage_0_output[2][8] ), .CP(clk), 
        .Q(\stage_0_retimer[2][8] ) );
  DFQD1 \stage_0_retimer_reg[2][7]  ( .D(\stage_0_output[2][7] ), .CP(clk), 
        .Q(\stage_0_retimer[2][7] ) );
  DFQD1 \stage_0_retimer_reg[2][6]  ( .D(\stage_0_output[2][6] ), .CP(clk), 
        .Q(\stage_0_retimer[2][6] ) );
  DFQD1 \stage_0_retimer_reg[2][5]  ( .D(\stage_0_output[2][5] ), .CP(clk), 
        .Q(\stage_0_retimer[2][5] ) );
  DFQD1 \stage_0_retimer_reg[2][4]  ( .D(\stage_0_output[2][4] ), .CP(clk), 
        .Q(\stage_0_retimer[2][4] ) );
  DFQD1 \stage_0_retimer_reg[2][3]  ( .D(\stage_0_output[2][3] ), .CP(clk), 
        .Q(\stage_0_retimer[2][3] ) );
  DFQD1 \stage_0_retimer_reg[2][2]  ( .D(\stage_0_output[2][2] ), .CP(clk), 
        .Q(\stage_0_retimer[2][2] ) );
  DFQD1 \stage_0_retimer_reg[2][1]  ( .D(\stage_0_output[2][1] ), .CP(clk), 
        .Q(\stage_0_retimer[2][1] ) );
  DFQD1 \stage_0_retimer_reg[2][0]  ( .D(\stage_0_output[2][0] ), .CP(clk), 
        .Q(\stage_0_retimer[2][0] ) );
  DFQD1 \stage_0_retimer_reg[1][19]  ( .D(\stage_0_output[1][19] ), .CP(clk), 
        .Q(\stage_0_retimer[1][19] ) );
  DFQD1 \stage_0_retimer_reg[1][18]  ( .D(\stage_0_output[1][18] ), .CP(clk), 
        .Q(\stage_0_retimer[1][18] ) );
  DFQD1 \stage_0_retimer_reg[1][17]  ( .D(\stage_0_output[1][17] ), .CP(clk), 
        .Q(\stage_0_retimer[1][17] ) );
  DFQD1 \stage_0_retimer_reg[1][16]  ( .D(\stage_0_output[1][16] ), .CP(clk), 
        .Q(\stage_0_retimer[1][16] ) );
  DFQD1 \stage_0_retimer_reg[1][15]  ( .D(\stage_0_output[1][15] ), .CP(clk), 
        .Q(\stage_0_retimer[1][15] ) );
  DFQD1 \stage_0_retimer_reg[1][14]  ( .D(\stage_0_output[1][14] ), .CP(clk), 
        .Q(\stage_0_retimer[1][14] ) );
  DFQD1 \stage_0_retimer_reg[1][13]  ( .D(\stage_0_output[1][13] ), .CP(clk), 
        .Q(\stage_0_retimer[1][13] ) );
  DFQD1 \stage_0_retimer_reg[1][12]  ( .D(\stage_0_output[1][12] ), .CP(clk), 
        .Q(\stage_0_retimer[1][12] ) );
  DFQD1 \stage_0_retimer_reg[1][11]  ( .D(\stage_0_output[1][11] ), .CP(clk), 
        .Q(\stage_0_retimer[1][11] ) );
  DFQD1 \stage_0_retimer_reg[1][10]  ( .D(\stage_0_output[1][10] ), .CP(clk), 
        .Q(\stage_0_retimer[1][10] ) );
  DFQD1 \stage_0_retimer_reg[1][9]  ( .D(\stage_0_output[1][9] ), .CP(clk), 
        .Q(\stage_0_retimer[1][9] ) );
  DFQD1 \stage_0_retimer_reg[1][8]  ( .D(\stage_0_output[1][8] ), .CP(clk), 
        .Q(\stage_0_retimer[1][8] ) );
  DFQD1 \stage_0_retimer_reg[1][7]  ( .D(\stage_0_output[1][7] ), .CP(clk), 
        .Q(\stage_0_retimer[1][7] ) );
  DFQD1 \stage_0_retimer_reg[1][6]  ( .D(\stage_0_output[1][6] ), .CP(clk), 
        .Q(\stage_0_retimer[1][6] ) );
  DFQD1 \stage_0_retimer_reg[1][5]  ( .D(\stage_0_output[1][5] ), .CP(clk), 
        .Q(\stage_0_retimer[1][5] ) );
  DFQD1 \stage_0_retimer_reg[1][4]  ( .D(\stage_0_output[1][4] ), .CP(clk), 
        .Q(\stage_0_retimer[1][4] ) );
  DFQD1 \stage_0_retimer_reg[1][3]  ( .D(\stage_0_output[1][3] ), .CP(clk), 
        .Q(\stage_0_retimer[1][3] ) );
  DFQD1 \stage_0_retimer_reg[1][2]  ( .D(\stage_0_output[1][2] ), .CP(clk), 
        .Q(\stage_0_retimer[1][2] ) );
  DFQD1 \stage_0_retimer_reg[1][1]  ( .D(\stage_0_output[1][1] ), .CP(clk), 
        .Q(\stage_0_retimer[1][1] ) );
  DFQD1 \stage_0_retimer_reg[1][0]  ( .D(\stage_0_output[1][0] ), .CP(clk), 
        .Q(\stage_0_retimer[1][0] ) );
  DFQD1 \stage_0_retimer_reg[0][19]  ( .D(\stage_0_output[0][19] ), .CP(clk), 
        .Q(\stage_0_retimer[0][19] ) );
  DFQD1 \stage_0_retimer_reg[0][18]  ( .D(\stage_0_output[0][18] ), .CP(clk), 
        .Q(\stage_0_retimer[0][18] ) );
  DFQD1 \stage_0_retimer_reg[0][17]  ( .D(\stage_0_output[0][17] ), .CP(clk), 
        .Q(\stage_0_retimer[0][17] ) );
  DFQD1 \stage_0_retimer_reg[0][16]  ( .D(\stage_0_output[0][16] ), .CP(clk), 
        .Q(\stage_0_retimer[0][16] ) );
  DFQD1 \stage_0_retimer_reg[0][15]  ( .D(\stage_0_output[0][15] ), .CP(clk), 
        .Q(\stage_0_retimer[0][15] ) );
  DFQD1 \stage_0_retimer_reg[0][14]  ( .D(\stage_0_output[0][14] ), .CP(clk), 
        .Q(\stage_0_retimer[0][14] ) );
  DFQD1 \stage_0_retimer_reg[0][13]  ( .D(\stage_0_output[0][13] ), .CP(clk), 
        .Q(\stage_0_retimer[0][13] ) );
  DFQD1 \stage_0_retimer_reg[0][12]  ( .D(\stage_0_output[0][12] ), .CP(clk), 
        .Q(\stage_0_retimer[0][12] ) );
  DFQD1 \stage_0_retimer_reg[0][11]  ( .D(\stage_0_output[0][11] ), .CP(clk), 
        .Q(\stage_0_retimer[0][11] ) );
  DFQD1 \stage_0_retimer_reg[0][10]  ( .D(\stage_0_output[0][10] ), .CP(clk), 
        .Q(\stage_0_retimer[0][10] ) );
  DFQD1 \stage_0_retimer_reg[0][9]  ( .D(\stage_0_output[0][9] ), .CP(clk), 
        .Q(\stage_0_retimer[0][9] ) );
  DFQD1 \stage_0_retimer_reg[0][8]  ( .D(\stage_0_output[0][8] ), .CP(clk), 
        .Q(\stage_0_retimer[0][8] ) );
  DFQD1 \stage_0_retimer_reg[0][7]  ( .D(\stage_0_output[0][7] ), .CP(clk), 
        .Q(\stage_0_retimer[0][7] ) );
  DFQD1 \stage_0_retimer_reg[0][6]  ( .D(\stage_0_output[0][6] ), .CP(clk), 
        .Q(\stage_0_retimer[0][6] ) );
  DFQD1 \stage_0_retimer_reg[0][5]  ( .D(\stage_0_output[0][5] ), .CP(clk), 
        .Q(\stage_0_retimer[0][5] ) );
  DFQD1 \stage_0_retimer_reg[0][4]  ( .D(\stage_0_output[0][4] ), .CP(clk), 
        .Q(\stage_0_retimer[0][4] ) );
  DFQD1 \stage_0_retimer_reg[0][3]  ( .D(\stage_0_output[0][3] ), .CP(clk), 
        .Q(\stage_0_retimer[0][3] ) );
  DFQD1 \stage_0_retimer_reg[0][2]  ( .D(\stage_0_output[0][2] ), .CP(clk), 
        .Q(\stage_0_retimer[0][2] ) );
  DFQD1 \stage_0_retimer_reg[0][1]  ( .D(\stage_0_output[0][1] ), .CP(clk), 
        .Q(\stage_0_retimer[0][1] ) );
  DFQD1 \stage_0_retimer_reg[0][0]  ( .D(\stage_0_output[0][0] ), .CP(clk), 
        .Q(\stage_0_retimer[0][0] ) );
  DFQD1 \stage_1_retimer_reg[7][19]  ( .D(\stage_1_output[7][19] ), .CP(clk), 
        .Q(\stage_1_retimer[7][19] ) );
  DFQD1 \stage_1_retimer_reg[7][18]  ( .D(\stage_1_output[7][18] ), .CP(clk), 
        .Q(\stage_1_retimer[7][18] ) );
  DFQD1 \stage_1_retimer_reg[7][17]  ( .D(\stage_1_output[7][17] ), .CP(clk), 
        .Q(\stage_1_retimer[7][17] ) );
  DFQD1 \stage_1_retimer_reg[7][16]  ( .D(\stage_1_output[7][16] ), .CP(clk), 
        .Q(\stage_1_retimer[7][16] ) );
  DFQD1 \stage_1_retimer_reg[7][15]  ( .D(\stage_1_output[7][15] ), .CP(clk), 
        .Q(\stage_1_retimer[7][15] ) );
  DFQD1 \stage_1_retimer_reg[7][14]  ( .D(\stage_1_output[7][14] ), .CP(clk), 
        .Q(\stage_1_retimer[7][14] ) );
  DFQD1 \stage_1_retimer_reg[7][13]  ( .D(\stage_1_output[7][13] ), .CP(clk), 
        .Q(\stage_1_retimer[7][13] ) );
  DFQD1 \stage_1_retimer_reg[7][12]  ( .D(\stage_1_output[7][12] ), .CP(clk), 
        .Q(\stage_1_retimer[7][12] ) );
  DFQD1 \stage_1_retimer_reg[7][11]  ( .D(\stage_1_output[7][11] ), .CP(clk), 
        .Q(\stage_1_retimer[7][11] ) );
  DFQD1 \stage_1_retimer_reg[7][10]  ( .D(\stage_1_output[7][10] ), .CP(clk), 
        .Q(\stage_1_retimer[7][10] ) );
  DFQD1 \stage_1_retimer_reg[7][9]  ( .D(\stage_1_output[7][9] ), .CP(clk), 
        .Q(\stage_1_retimer[7][9] ) );
  DFQD1 \stage_1_retimer_reg[7][8]  ( .D(\stage_1_output[7][8] ), .CP(clk), 
        .Q(\stage_1_retimer[7][8] ) );
  DFQD1 \stage_1_retimer_reg[7][7]  ( .D(\stage_1_output[7][7] ), .CP(clk), 
        .Q(\stage_1_retimer[7][7] ) );
  DFQD1 \stage_1_retimer_reg[7][6]  ( .D(\stage_1_output[7][6] ), .CP(clk), 
        .Q(\stage_1_retimer[7][6] ) );
  DFQD1 \stage_1_retimer_reg[7][5]  ( .D(\stage_1_output[7][5] ), .CP(clk), 
        .Q(\stage_1_retimer[7][5] ) );
  DFQD1 \stage_1_retimer_reg[7][4]  ( .D(\stage_1_output[7][4] ), .CP(clk), 
        .Q(\stage_1_retimer[7][4] ) );
  DFQD1 \stage_1_retimer_reg[7][3]  ( .D(\stage_1_output[7][3] ), .CP(clk), 
        .Q(\stage_1_retimer[7][3] ) );
  DFQD1 \stage_1_retimer_reg[7][2]  ( .D(\stage_1_output[7][2] ), .CP(clk), 
        .Q(\stage_1_retimer[7][2] ) );
  DFQD1 \stage_1_retimer_reg[7][1]  ( .D(\stage_1_output[7][1] ), .CP(clk), 
        .Q(\stage_1_retimer[7][1] ) );
  DFQD1 \stage_1_retimer_reg[7][0]  ( .D(\stage_1_output[7][0] ), .CP(clk), 
        .Q(\stage_1_retimer[7][0] ) );
  DFQD1 \stage_1_retimer_reg[6][19]  ( .D(\stage_1_output[6][19] ), .CP(clk), 
        .Q(\stage_1_retimer[6][19] ) );
  DFQD1 \stage_1_retimer_reg[6][18]  ( .D(\stage_1_output[6][18] ), .CP(clk), 
        .Q(\stage_1_retimer[6][18] ) );
  DFQD1 \stage_1_retimer_reg[6][17]  ( .D(\stage_1_output[6][17] ), .CP(clk), 
        .Q(\stage_1_retimer[6][17] ) );
  DFQD1 \stage_1_retimer_reg[6][16]  ( .D(\stage_1_output[6][16] ), .CP(clk), 
        .Q(\stage_1_retimer[6][16] ) );
  DFQD1 \stage_1_retimer_reg[6][15]  ( .D(\stage_1_output[6][15] ), .CP(clk), 
        .Q(\stage_1_retimer[6][15] ) );
  DFQD1 \stage_1_retimer_reg[6][14]  ( .D(\stage_1_output[6][14] ), .CP(clk), 
        .Q(\stage_1_retimer[6][14] ) );
  DFQD1 \stage_1_retimer_reg[6][13]  ( .D(\stage_1_output[6][13] ), .CP(clk), 
        .Q(\stage_1_retimer[6][13] ) );
  DFQD1 \stage_1_retimer_reg[6][12]  ( .D(\stage_1_output[6][12] ), .CP(clk), 
        .Q(\stage_1_retimer[6][12] ) );
  DFQD1 \stage_1_retimer_reg[6][11]  ( .D(\stage_1_output[6][11] ), .CP(clk), 
        .Q(\stage_1_retimer[6][11] ) );
  DFQD1 \stage_1_retimer_reg[6][10]  ( .D(\stage_1_output[6][10] ), .CP(clk), 
        .Q(\stage_1_retimer[6][10] ) );
  DFQD1 \stage_1_retimer_reg[6][9]  ( .D(\stage_1_output[6][9] ), .CP(clk), 
        .Q(\stage_1_retimer[6][9] ) );
  DFQD1 \stage_1_retimer_reg[6][8]  ( .D(\stage_1_output[6][8] ), .CP(clk), 
        .Q(\stage_1_retimer[6][8] ) );
  DFQD1 \stage_1_retimer_reg[6][7]  ( .D(\stage_1_output[6][7] ), .CP(clk), 
        .Q(\stage_1_retimer[6][7] ) );
  DFQD1 \stage_1_retimer_reg[6][6]  ( .D(\stage_1_output[6][6] ), .CP(clk), 
        .Q(\stage_1_retimer[6][6] ) );
  DFQD1 \stage_1_retimer_reg[6][5]  ( .D(\stage_1_output[6][5] ), .CP(clk), 
        .Q(\stage_1_retimer[6][5] ) );
  DFQD1 \stage_1_retimer_reg[6][4]  ( .D(\stage_1_output[6][4] ), .CP(clk), 
        .Q(\stage_1_retimer[6][4] ) );
  DFQD1 \stage_1_retimer_reg[6][3]  ( .D(\stage_1_output[6][3] ), .CP(clk), 
        .Q(\stage_1_retimer[6][3] ) );
  DFQD1 \stage_1_retimer_reg[6][2]  ( .D(\stage_1_output[6][2] ), .CP(clk), 
        .Q(\stage_1_retimer[6][2] ) );
  DFQD1 \stage_1_retimer_reg[6][1]  ( .D(\stage_1_output[6][1] ), .CP(clk), 
        .Q(\stage_1_retimer[6][1] ) );
  DFQD1 \stage_1_retimer_reg[6][0]  ( .D(\stage_1_output[6][0] ), .CP(clk), 
        .Q(\stage_1_retimer[6][0] ) );
  DFQD1 \stage_1_retimer_reg[5][19]  ( .D(\stage_1_output[5][19] ), .CP(clk), 
        .Q(\stage_1_retimer[5][19] ) );
  DFQD1 \stage_1_retimer_reg[5][18]  ( .D(\stage_1_output[5][18] ), .CP(clk), 
        .Q(\stage_1_retimer[5][18] ) );
  DFQD1 \stage_1_retimer_reg[5][17]  ( .D(\stage_1_output[5][17] ), .CP(clk), 
        .Q(\stage_1_retimer[5][17] ) );
  DFQD1 \stage_1_retimer_reg[5][16]  ( .D(\stage_1_output[5][16] ), .CP(clk), 
        .Q(\stage_1_retimer[5][16] ) );
  DFQD1 \stage_1_retimer_reg[5][15]  ( .D(\stage_1_output[5][15] ), .CP(clk), 
        .Q(\stage_1_retimer[5][15] ) );
  DFQD1 \stage_1_retimer_reg[5][14]  ( .D(\stage_1_output[5][14] ), .CP(clk), 
        .Q(\stage_1_retimer[5][14] ) );
  DFQD1 \stage_1_retimer_reg[5][13]  ( .D(\stage_1_output[5][13] ), .CP(clk), 
        .Q(\stage_1_retimer[5][13] ) );
  DFQD1 \stage_1_retimer_reg[5][12]  ( .D(\stage_1_output[5][12] ), .CP(clk), 
        .Q(\stage_1_retimer[5][12] ) );
  DFQD1 \stage_1_retimer_reg[5][11]  ( .D(\stage_1_output[5][11] ), .CP(clk), 
        .Q(\stage_1_retimer[5][11] ) );
  DFQD1 \stage_1_retimer_reg[5][10]  ( .D(\stage_1_output[5][10] ), .CP(clk), 
        .Q(\stage_1_retimer[5][10] ) );
  DFQD1 \stage_1_retimer_reg[5][9]  ( .D(\stage_1_output[5][9] ), .CP(clk), 
        .Q(\stage_1_retimer[5][9] ) );
  DFQD1 \stage_1_retimer_reg[5][8]  ( .D(\stage_1_output[5][8] ), .CP(clk), 
        .Q(\stage_1_retimer[5][8] ) );
  DFQD1 \stage_1_retimer_reg[5][7]  ( .D(\stage_1_output[5][7] ), .CP(clk), 
        .Q(\stage_1_retimer[5][7] ) );
  DFQD1 \stage_1_retimer_reg[5][6]  ( .D(\stage_1_output[5][6] ), .CP(clk), 
        .Q(\stage_1_retimer[5][6] ) );
  DFQD1 \stage_1_retimer_reg[5][5]  ( .D(\stage_1_output[5][5] ), .CP(clk), 
        .Q(\stage_1_retimer[5][5] ) );
  DFQD1 \stage_1_retimer_reg[5][4]  ( .D(\stage_1_output[5][4] ), .CP(clk), 
        .Q(\stage_1_retimer[5][4] ) );
  DFQD1 \stage_1_retimer_reg[5][3]  ( .D(\stage_1_output[5][3] ), .CP(clk), 
        .Q(\stage_1_retimer[5][3] ) );
  DFQD1 \stage_1_retimer_reg[5][2]  ( .D(\stage_1_output[5][2] ), .CP(clk), 
        .Q(\stage_1_retimer[5][2] ) );
  DFQD1 \stage_1_retimer_reg[5][1]  ( .D(\stage_1_output[5][1] ), .CP(clk), 
        .Q(\stage_1_retimer[5][1] ) );
  DFQD1 \stage_1_retimer_reg[5][0]  ( .D(\stage_1_output[5][0] ), .CP(clk), 
        .Q(\stage_1_retimer[5][0] ) );
  DFQD1 \stage_1_retimer_reg[4][19]  ( .D(\stage_1_output[4][19] ), .CP(clk), 
        .Q(\stage_1_retimer[4][19] ) );
  DFQD1 \stage_1_retimer_reg[4][18]  ( .D(\stage_1_output[4][18] ), .CP(clk), 
        .Q(\stage_1_retimer[4][18] ) );
  DFQD1 \stage_1_retimer_reg[4][17]  ( .D(\stage_1_output[4][17] ), .CP(clk), 
        .Q(\stage_1_retimer[4][17] ) );
  DFQD1 \stage_1_retimer_reg[4][16]  ( .D(\stage_1_output[4][16] ), .CP(clk), 
        .Q(\stage_1_retimer[4][16] ) );
  DFQD1 \stage_1_retimer_reg[4][15]  ( .D(\stage_1_output[4][15] ), .CP(clk), 
        .Q(\stage_1_retimer[4][15] ) );
  DFQD1 \stage_1_retimer_reg[4][14]  ( .D(\stage_1_output[4][14] ), .CP(clk), 
        .Q(\stage_1_retimer[4][14] ) );
  DFQD1 \stage_1_retimer_reg[4][13]  ( .D(\stage_1_output[4][13] ), .CP(clk), 
        .Q(\stage_1_retimer[4][13] ) );
  DFQD1 \stage_1_retimer_reg[4][12]  ( .D(\stage_1_output[4][12] ), .CP(clk), 
        .Q(\stage_1_retimer[4][12] ) );
  DFQD1 \stage_1_retimer_reg[4][11]  ( .D(\stage_1_output[4][11] ), .CP(clk), 
        .Q(\stage_1_retimer[4][11] ) );
  DFQD1 \stage_1_retimer_reg[4][10]  ( .D(\stage_1_output[4][10] ), .CP(clk), 
        .Q(\stage_1_retimer[4][10] ) );
  DFQD1 \stage_1_retimer_reg[4][9]  ( .D(\stage_1_output[4][9] ), .CP(clk), 
        .Q(\stage_1_retimer[4][9] ) );
  DFQD1 \stage_1_retimer_reg[4][8]  ( .D(\stage_1_output[4][8] ), .CP(clk), 
        .Q(\stage_1_retimer[4][8] ) );
  DFQD1 \stage_1_retimer_reg[4][7]  ( .D(\stage_1_output[4][7] ), .CP(clk), 
        .Q(\stage_1_retimer[4][7] ) );
  DFQD1 \stage_1_retimer_reg[4][6]  ( .D(\stage_1_output[4][6] ), .CP(clk), 
        .Q(\stage_1_retimer[4][6] ) );
  DFQD1 \stage_1_retimer_reg[4][5]  ( .D(\stage_1_output[4][5] ), .CP(clk), 
        .Q(\stage_1_retimer[4][5] ) );
  DFQD1 \stage_1_retimer_reg[4][4]  ( .D(\stage_1_output[4][4] ), .CP(clk), 
        .Q(\stage_1_retimer[4][4] ) );
  DFQD1 \stage_1_retimer_reg[4][3]  ( .D(\stage_1_output[4][3] ), .CP(clk), 
        .Q(\stage_1_retimer[4][3] ) );
  DFQD1 \stage_1_retimer_reg[4][2]  ( .D(\stage_1_output[4][2] ), .CP(clk), 
        .Q(\stage_1_retimer[4][2] ) );
  DFQD1 \stage_1_retimer_reg[4][1]  ( .D(\stage_1_output[4][1] ), .CP(clk), 
        .Q(\stage_1_retimer[4][1] ) );
  DFQD1 \stage_1_retimer_reg[4][0]  ( .D(\stage_1_output[4][0] ), .CP(clk), 
        .Q(\stage_1_retimer[4][0] ) );
  DFQD1 \stage_1_retimer_reg[3][19]  ( .D(\stage_1_output[3][19] ), .CP(clk), 
        .Q(\stage_1_retimer[3][19] ) );
  DFQD1 \stage_1_retimer_reg[3][18]  ( .D(\stage_1_output[3][18] ), .CP(clk), 
        .Q(\stage_1_retimer[3][18] ) );
  DFQD1 \stage_1_retimer_reg[3][17]  ( .D(\stage_1_output[3][17] ), .CP(clk), 
        .Q(\stage_1_retimer[3][17] ) );
  DFQD1 \stage_1_retimer_reg[3][16]  ( .D(\stage_1_output[3][16] ), .CP(clk), 
        .Q(\stage_1_retimer[3][16] ) );
  DFQD1 \stage_1_retimer_reg[3][15]  ( .D(\stage_1_output[3][15] ), .CP(clk), 
        .Q(\stage_1_retimer[3][15] ) );
  DFQD1 \stage_1_retimer_reg[3][14]  ( .D(\stage_1_output[3][14] ), .CP(clk), 
        .Q(\stage_1_retimer[3][14] ) );
  DFQD1 \stage_1_retimer_reg[3][13]  ( .D(\stage_1_output[3][13] ), .CP(clk), 
        .Q(\stage_1_retimer[3][13] ) );
  DFQD1 \stage_1_retimer_reg[3][12]  ( .D(\stage_1_output[3][12] ), .CP(clk), 
        .Q(\stage_1_retimer[3][12] ) );
  DFQD1 \stage_1_retimer_reg[3][11]  ( .D(\stage_1_output[3][11] ), .CP(clk), 
        .Q(\stage_1_retimer[3][11] ) );
  DFQD1 \stage_1_retimer_reg[3][10]  ( .D(\stage_1_output[3][10] ), .CP(clk), 
        .Q(\stage_1_retimer[3][10] ) );
  DFQD1 \stage_1_retimer_reg[3][9]  ( .D(\stage_1_output[3][9] ), .CP(clk), 
        .Q(\stage_1_retimer[3][9] ) );
  DFQD1 \stage_1_retimer_reg[3][8]  ( .D(\stage_1_output[3][8] ), .CP(clk), 
        .Q(\stage_1_retimer[3][8] ) );
  DFQD1 \stage_1_retimer_reg[3][7]  ( .D(\stage_1_output[3][7] ), .CP(clk), 
        .Q(\stage_1_retimer[3][7] ) );
  DFQD1 \stage_1_retimer_reg[3][6]  ( .D(\stage_1_output[3][6] ), .CP(clk), 
        .Q(\stage_1_retimer[3][6] ) );
  DFQD1 \stage_1_retimer_reg[3][5]  ( .D(\stage_1_output[3][5] ), .CP(clk), 
        .Q(\stage_1_retimer[3][5] ) );
  DFQD1 \stage_1_retimer_reg[3][4]  ( .D(\stage_1_output[3][4] ), .CP(clk), 
        .Q(\stage_1_retimer[3][4] ) );
  DFQD1 \stage_1_retimer_reg[3][3]  ( .D(\stage_1_output[3][3] ), .CP(clk), 
        .Q(\stage_1_retimer[3][3] ) );
  DFQD1 \stage_1_retimer_reg[3][2]  ( .D(\stage_1_output[3][2] ), .CP(clk), 
        .Q(\stage_1_retimer[3][2] ) );
  DFQD1 \stage_1_retimer_reg[3][1]  ( .D(\stage_1_output[3][1] ), .CP(clk), 
        .Q(\stage_1_retimer[3][1] ) );
  DFQD1 \stage_1_retimer_reg[3][0]  ( .D(\stage_1_output[3][0] ), .CP(clk), 
        .Q(\stage_1_retimer[3][0] ) );
  DFQD1 \stage_1_retimer_reg[2][19]  ( .D(\stage_1_output[2][19] ), .CP(clk), 
        .Q(\stage_1_retimer[2][19] ) );
  DFQD1 \stage_1_retimer_reg[2][18]  ( .D(\stage_1_output[2][18] ), .CP(clk), 
        .Q(\stage_1_retimer[2][18] ) );
  DFQD1 \stage_1_retimer_reg[2][17]  ( .D(\stage_1_output[2][17] ), .CP(clk), 
        .Q(\stage_1_retimer[2][17] ) );
  DFQD1 \stage_1_retimer_reg[2][16]  ( .D(\stage_1_output[2][16] ), .CP(clk), 
        .Q(\stage_1_retimer[2][16] ) );
  DFQD1 \stage_1_retimer_reg[2][15]  ( .D(\stage_1_output[2][15] ), .CP(clk), 
        .Q(\stage_1_retimer[2][15] ) );
  DFQD1 \stage_1_retimer_reg[2][14]  ( .D(\stage_1_output[2][14] ), .CP(clk), 
        .Q(\stage_1_retimer[2][14] ) );
  DFQD1 \stage_1_retimer_reg[2][13]  ( .D(\stage_1_output[2][13] ), .CP(clk), 
        .Q(\stage_1_retimer[2][13] ) );
  DFQD1 \stage_1_retimer_reg[2][12]  ( .D(\stage_1_output[2][12] ), .CP(clk), 
        .Q(\stage_1_retimer[2][12] ) );
  DFQD1 \stage_1_retimer_reg[2][11]  ( .D(\stage_1_output[2][11] ), .CP(clk), 
        .Q(\stage_1_retimer[2][11] ) );
  DFQD1 \stage_1_retimer_reg[2][10]  ( .D(\stage_1_output[2][10] ), .CP(clk), 
        .Q(\stage_1_retimer[2][10] ) );
  DFQD1 \stage_1_retimer_reg[2][9]  ( .D(\stage_1_output[2][9] ), .CP(clk), 
        .Q(\stage_1_retimer[2][9] ) );
  DFQD1 \stage_1_retimer_reg[2][8]  ( .D(\stage_1_output[2][8] ), .CP(clk), 
        .Q(\stage_1_retimer[2][8] ) );
  DFQD1 \stage_1_retimer_reg[2][7]  ( .D(\stage_1_output[2][7] ), .CP(clk), 
        .Q(\stage_1_retimer[2][7] ) );
  DFQD1 \stage_1_retimer_reg[2][6]  ( .D(\stage_1_output[2][6] ), .CP(clk), 
        .Q(\stage_1_retimer[2][6] ) );
  DFQD1 \stage_1_retimer_reg[2][5]  ( .D(\stage_1_output[2][5] ), .CP(clk), 
        .Q(\stage_1_retimer[2][5] ) );
  DFQD1 \stage_1_retimer_reg[2][4]  ( .D(\stage_1_output[2][4] ), .CP(clk), 
        .Q(\stage_1_retimer[2][4] ) );
  DFQD1 \stage_1_retimer_reg[2][3]  ( .D(\stage_1_output[2][3] ), .CP(clk), 
        .Q(\stage_1_retimer[2][3] ) );
  DFQD1 \stage_1_retimer_reg[2][2]  ( .D(\stage_1_output[2][2] ), .CP(clk), 
        .Q(\stage_1_retimer[2][2] ) );
  DFQD1 \stage_1_retimer_reg[2][1]  ( .D(\stage_1_output[2][1] ), .CP(clk), 
        .Q(\stage_1_retimer[2][1] ) );
  DFQD1 \stage_1_retimer_reg[2][0]  ( .D(\stage_1_output[2][0] ), .CP(clk), 
        .Q(\stage_1_retimer[2][0] ) );
  DFQD1 \stage_1_retimer_reg[1][19]  ( .D(\stage_1_output[1][19] ), .CP(clk), 
        .Q(\stage_1_retimer[1][19] ) );
  DFQD1 \stage_1_retimer_reg[1][18]  ( .D(\stage_1_output[1][18] ), .CP(clk), 
        .Q(\stage_1_retimer[1][18] ) );
  DFQD1 \stage_1_retimer_reg[1][17]  ( .D(\stage_1_output[1][17] ), .CP(clk), 
        .Q(\stage_1_retimer[1][17] ) );
  DFQD1 \stage_1_retimer_reg[1][16]  ( .D(\stage_1_output[1][16] ), .CP(clk), 
        .Q(\stage_1_retimer[1][16] ) );
  DFQD1 \stage_1_retimer_reg[1][15]  ( .D(\stage_1_output[1][15] ), .CP(clk), 
        .Q(\stage_1_retimer[1][15] ) );
  DFQD1 \stage_1_retimer_reg[1][14]  ( .D(\stage_1_output[1][14] ), .CP(clk), 
        .Q(\stage_1_retimer[1][14] ) );
  DFQD1 \stage_1_retimer_reg[1][13]  ( .D(\stage_1_output[1][13] ), .CP(clk), 
        .Q(\stage_1_retimer[1][13] ) );
  DFQD1 \stage_1_retimer_reg[1][12]  ( .D(\stage_1_output[1][12] ), .CP(clk), 
        .Q(\stage_1_retimer[1][12] ) );
  DFQD1 \stage_1_retimer_reg[1][11]  ( .D(\stage_1_output[1][11] ), .CP(clk), 
        .Q(\stage_1_retimer[1][11] ) );
  DFQD1 \stage_1_retimer_reg[1][10]  ( .D(\stage_1_output[1][10] ), .CP(clk), 
        .Q(\stage_1_retimer[1][10] ) );
  DFQD1 \stage_1_retimer_reg[1][9]  ( .D(\stage_1_output[1][9] ), .CP(clk), 
        .Q(\stage_1_retimer[1][9] ) );
  DFQD1 \stage_1_retimer_reg[1][8]  ( .D(\stage_1_output[1][8] ), .CP(clk), 
        .Q(\stage_1_retimer[1][8] ) );
  DFQD1 \stage_1_retimer_reg[1][7]  ( .D(\stage_1_output[1][7] ), .CP(clk), 
        .Q(\stage_1_retimer[1][7] ) );
  DFQD1 \stage_1_retimer_reg[1][6]  ( .D(\stage_1_output[1][6] ), .CP(clk), 
        .Q(\stage_1_retimer[1][6] ) );
  DFQD1 \stage_1_retimer_reg[1][5]  ( .D(\stage_1_output[1][5] ), .CP(clk), 
        .Q(\stage_1_retimer[1][5] ) );
  DFQD1 \stage_1_retimer_reg[1][4]  ( .D(\stage_1_output[1][4] ), .CP(clk), 
        .Q(\stage_1_retimer[1][4] ) );
  DFQD1 \stage_1_retimer_reg[1][3]  ( .D(\stage_1_output[1][3] ), .CP(clk), 
        .Q(\stage_1_retimer[1][3] ) );
  DFQD1 \stage_1_retimer_reg[1][2]  ( .D(\stage_1_output[1][2] ), .CP(clk), 
        .Q(\stage_1_retimer[1][2] ) );
  DFQD1 \stage_1_retimer_reg[1][1]  ( .D(\stage_1_output[1][1] ), .CP(clk), 
        .Q(\stage_1_retimer[1][1] ) );
  DFQD1 \stage_1_retimer_reg[1][0]  ( .D(\stage_1_output[1][0] ), .CP(clk), 
        .Q(\stage_1_retimer[1][0] ) );
  DFQD1 \stage_1_retimer_reg[0][19]  ( .D(\stage_1_output[0][19] ), .CP(clk), 
        .Q(\stage_1_retimer[0][19] ) );
  DFQD1 \stage_1_retimer_reg[0][18]  ( .D(\stage_1_output[0][18] ), .CP(clk), 
        .Q(\stage_1_retimer[0][18] ) );
  DFQD1 \stage_1_retimer_reg[0][17]  ( .D(\stage_1_output[0][17] ), .CP(clk), 
        .Q(\stage_1_retimer[0][17] ) );
  DFQD1 \stage_1_retimer_reg[0][16]  ( .D(\stage_1_output[0][16] ), .CP(clk), 
        .Q(\stage_1_retimer[0][16] ) );
  DFQD1 \stage_1_retimer_reg[0][15]  ( .D(\stage_1_output[0][15] ), .CP(clk), 
        .Q(\stage_1_retimer[0][15] ) );
  DFQD1 \stage_1_retimer_reg[0][14]  ( .D(\stage_1_output[0][14] ), .CP(clk), 
        .Q(\stage_1_retimer[0][14] ) );
  DFQD1 \stage_1_retimer_reg[0][13]  ( .D(\stage_1_output[0][13] ), .CP(clk), 
        .Q(\stage_1_retimer[0][13] ) );
  DFQD1 \stage_1_retimer_reg[0][12]  ( .D(\stage_1_output[0][12] ), .CP(clk), 
        .Q(\stage_1_retimer[0][12] ) );
  DFQD1 \stage_1_retimer_reg[0][11]  ( .D(\stage_1_output[0][11] ), .CP(clk), 
        .Q(\stage_1_retimer[0][11] ) );
  DFQD1 \stage_1_retimer_reg[0][10]  ( .D(\stage_1_output[0][10] ), .CP(clk), 
        .Q(\stage_1_retimer[0][10] ) );
  DFQD1 \stage_1_retimer_reg[0][9]  ( .D(\stage_1_output[0][9] ), .CP(clk), 
        .Q(\stage_1_retimer[0][9] ) );
  DFQD1 \stage_1_retimer_reg[0][8]  ( .D(\stage_1_output[0][8] ), .CP(clk), 
        .Q(\stage_1_retimer[0][8] ) );
  DFQD1 \stage_1_retimer_reg[0][7]  ( .D(\stage_1_output[0][7] ), .CP(clk), 
        .Q(\stage_1_retimer[0][7] ) );
  DFQD1 \stage_1_retimer_reg[0][6]  ( .D(\stage_1_output[0][6] ), .CP(clk), 
        .Q(\stage_1_retimer[0][6] ) );
  DFQD1 \stage_1_retimer_reg[0][5]  ( .D(\stage_1_output[0][5] ), .CP(clk), 
        .Q(\stage_1_retimer[0][5] ) );
  DFQD1 \stage_1_retimer_reg[0][4]  ( .D(\stage_1_output[0][4] ), .CP(clk), 
        .Q(\stage_1_retimer[0][4] ) );
  DFQD1 \stage_1_retimer_reg[0][3]  ( .D(\stage_1_output[0][3] ), .CP(clk), 
        .Q(\stage_1_retimer[0][3] ) );
  DFQD1 \stage_1_retimer_reg[0][2]  ( .D(\stage_1_output[0][2] ), .CP(clk), 
        .Q(\stage_1_retimer[0][2] ) );
  DFQD1 \stage_1_retimer_reg[0][1]  ( .D(\stage_1_output[0][1] ), .CP(clk), 
        .Q(\stage_1_retimer[0][1] ) );
  DFQD1 \stage_1_retimer_reg[0][0]  ( .D(\stage_1_output[0][0] ), .CP(clk), 
        .Q(\stage_1_retimer[0][0] ) );
  DFQD1 \stage_2_retimer_reg[7][19]  ( .D(\stage_2_output[7][19] ), .CP(clk), 
        .Q(\stage_2_retimer[7][19] ) );
  DFQD1 \stage_2_retimer_reg[7][18]  ( .D(\stage_2_output[7][18] ), .CP(clk), 
        .Q(\stage_2_retimer[7][18] ) );
  DFQD1 \stage_2_retimer_reg[7][17]  ( .D(\stage_2_output[7][17] ), .CP(clk), 
        .Q(\stage_2_retimer[7][17] ) );
  DFQD1 \stage_2_retimer_reg[7][16]  ( .D(\stage_2_output[7][16] ), .CP(clk), 
        .Q(\stage_2_retimer[7][16] ) );
  DFQD1 \stage_2_retimer_reg[7][15]  ( .D(\stage_2_output[7][15] ), .CP(clk), 
        .Q(\stage_2_retimer[7][15] ) );
  DFQD1 \stage_2_retimer_reg[7][14]  ( .D(\stage_2_output[7][14] ), .CP(clk), 
        .Q(\stage_2_retimer[7][14] ) );
  DFQD1 \stage_2_retimer_reg[7][13]  ( .D(\stage_2_output[7][13] ), .CP(clk), 
        .Q(\stage_2_retimer[7][13] ) );
  DFQD1 \stage_2_retimer_reg[7][12]  ( .D(\stage_2_output[7][12] ), .CP(clk), 
        .Q(\stage_2_retimer[7][12] ) );
  DFQD1 \stage_2_retimer_reg[7][11]  ( .D(\stage_2_output[7][11] ), .CP(clk), 
        .Q(\stage_2_retimer[7][11] ) );
  DFQD1 \stage_2_retimer_reg[7][10]  ( .D(\stage_2_output[7][10] ), .CP(clk), 
        .Q(\stage_2_retimer[7][10] ) );
  DFQD1 \stage_2_retimer_reg[7][9]  ( .D(\stage_2_output[7][9] ), .CP(clk), 
        .Q(\stage_2_retimer[7][9] ) );
  DFQD1 \stage_2_retimer_reg[7][8]  ( .D(\stage_2_output[7][8] ), .CP(clk), 
        .Q(\stage_2_retimer[7][8] ) );
  DFQD1 \stage_2_retimer_reg[7][7]  ( .D(\stage_2_output[7][7] ), .CP(clk), 
        .Q(\stage_2_retimer[7][7] ) );
  DFQD1 \stage_2_retimer_reg[7][6]  ( .D(\stage_2_output[7][6] ), .CP(clk), 
        .Q(\stage_2_retimer[7][6] ) );
  DFQD1 \stage_2_retimer_reg[7][5]  ( .D(\stage_2_output[7][5] ), .CP(clk), 
        .Q(\stage_2_retimer[7][5] ) );
  DFQD1 \stage_2_retimer_reg[7][4]  ( .D(\stage_2_output[7][4] ), .CP(clk), 
        .Q(\stage_2_retimer[7][4] ) );
  DFQD1 \stage_2_retimer_reg[7][3]  ( .D(\stage_2_output[7][3] ), .CP(clk), 
        .Q(\stage_2_retimer[7][3] ) );
  DFQD1 \stage_2_retimer_reg[7][2]  ( .D(\stage_2_output[7][2] ), .CP(clk), 
        .Q(\stage_2_retimer[7][2] ) );
  DFQD1 \stage_2_retimer_reg[7][1]  ( .D(\stage_2_output[7][1] ), .CP(clk), 
        .Q(\stage_2_retimer[7][1] ) );
  DFQD1 \stage_2_retimer_reg[7][0]  ( .D(\stage_2_output[7][0] ), .CP(clk), 
        .Q(\stage_2_retimer[7][0] ) );
  DFQD1 \stage_2_retimer_reg[6][19]  ( .D(\stage_2_output[6][19] ), .CP(clk), 
        .Q(\stage_2_retimer[6][19] ) );
  DFQD1 \stage_2_retimer_reg[6][18]  ( .D(\stage_2_output[6][18] ), .CP(clk), 
        .Q(\stage_2_retimer[6][18] ) );
  DFQD1 \stage_2_retimer_reg[6][17]  ( .D(\stage_2_output[6][17] ), .CP(clk), 
        .Q(\stage_2_retimer[6][17] ) );
  DFQD1 \stage_2_retimer_reg[6][16]  ( .D(\stage_2_output[6][16] ), .CP(clk), 
        .Q(\stage_2_retimer[6][16] ) );
  DFQD1 \stage_2_retimer_reg[6][15]  ( .D(\stage_2_output[6][15] ), .CP(clk), 
        .Q(\stage_2_retimer[6][15] ) );
  DFQD1 \stage_2_retimer_reg[6][14]  ( .D(\stage_2_output[6][14] ), .CP(clk), 
        .Q(\stage_2_retimer[6][14] ) );
  DFQD1 \stage_2_retimer_reg[6][13]  ( .D(\stage_2_output[6][13] ), .CP(clk), 
        .Q(\stage_2_retimer[6][13] ) );
  DFQD1 \stage_2_retimer_reg[6][12]  ( .D(\stage_2_output[6][12] ), .CP(clk), 
        .Q(\stage_2_retimer[6][12] ) );
  DFQD1 \stage_2_retimer_reg[6][11]  ( .D(\stage_2_output[6][11] ), .CP(clk), 
        .Q(\stage_2_retimer[6][11] ) );
  DFQD1 \stage_2_retimer_reg[6][10]  ( .D(\stage_2_output[6][10] ), .CP(clk), 
        .Q(\stage_2_retimer[6][10] ) );
  DFQD1 \stage_2_retimer_reg[6][9]  ( .D(\stage_2_output[6][9] ), .CP(clk), 
        .Q(\stage_2_retimer[6][9] ) );
  DFQD1 \stage_2_retimer_reg[6][8]  ( .D(\stage_2_output[6][8] ), .CP(clk), 
        .Q(\stage_2_retimer[6][8] ) );
  DFQD1 \stage_2_retimer_reg[6][7]  ( .D(\stage_2_output[6][7] ), .CP(clk), 
        .Q(\stage_2_retimer[6][7] ) );
  DFQD1 \stage_2_retimer_reg[6][6]  ( .D(\stage_2_output[6][6] ), .CP(clk), 
        .Q(\stage_2_retimer[6][6] ) );
  DFQD1 \stage_2_retimer_reg[6][5]  ( .D(\stage_2_output[6][5] ), .CP(clk), 
        .Q(\stage_2_retimer[6][5] ) );
  DFQD1 \stage_2_retimer_reg[6][4]  ( .D(\stage_2_output[6][4] ), .CP(clk), 
        .Q(\stage_2_retimer[6][4] ) );
  DFQD1 \stage_2_retimer_reg[6][3]  ( .D(\stage_2_output[6][3] ), .CP(clk), 
        .Q(\stage_2_retimer[6][3] ) );
  DFQD1 \stage_2_retimer_reg[6][2]  ( .D(\stage_2_output[6][2] ), .CP(clk), 
        .Q(\stage_2_retimer[6][2] ) );
  DFQD1 \stage_2_retimer_reg[6][1]  ( .D(\stage_2_output[6][1] ), .CP(clk), 
        .Q(\stage_2_retimer[6][1] ) );
  DFQD1 \stage_2_retimer_reg[6][0]  ( .D(\stage_2_output[6][0] ), .CP(clk), 
        .Q(\stage_2_retimer[6][0] ) );
  DFQD1 \stage_2_retimer_reg[5][19]  ( .D(\stage_2_output[5][19] ), .CP(clk), 
        .Q(\stage_2_retimer[5][19] ) );
  DFQD1 \stage_2_retimer_reg[5][18]  ( .D(\stage_2_output[5][18] ), .CP(clk), 
        .Q(\stage_2_retimer[5][18] ) );
  DFQD1 \stage_2_retimer_reg[5][17]  ( .D(\stage_2_output[5][17] ), .CP(clk), 
        .Q(\stage_2_retimer[5][17] ) );
  DFQD1 \stage_2_retimer_reg[5][16]  ( .D(\stage_2_output[5][16] ), .CP(clk), 
        .Q(\stage_2_retimer[5][16] ) );
  DFQD1 \stage_2_retimer_reg[5][15]  ( .D(\stage_2_output[5][15] ), .CP(clk), 
        .Q(\stage_2_retimer[5][15] ) );
  DFQD1 \stage_2_retimer_reg[5][14]  ( .D(\stage_2_output[5][14] ), .CP(clk), 
        .Q(\stage_2_retimer[5][14] ) );
  DFQD1 \stage_2_retimer_reg[5][13]  ( .D(\stage_2_output[5][13] ), .CP(clk), 
        .Q(\stage_2_retimer[5][13] ) );
  DFQD1 \stage_2_retimer_reg[5][12]  ( .D(\stage_2_output[5][12] ), .CP(clk), 
        .Q(\stage_2_retimer[5][12] ) );
  DFQD1 \stage_2_retimer_reg[5][11]  ( .D(\stage_2_output[5][11] ), .CP(clk), 
        .Q(\stage_2_retimer[5][11] ) );
  DFQD1 \stage_2_retimer_reg[5][10]  ( .D(\stage_2_output[5][10] ), .CP(clk), 
        .Q(\stage_2_retimer[5][10] ) );
  DFQD1 \stage_2_retimer_reg[5][9]  ( .D(\stage_2_output[5][9] ), .CP(clk), 
        .Q(\stage_2_retimer[5][9] ) );
  DFQD1 \stage_2_retimer_reg[5][8]  ( .D(\stage_2_output[5][8] ), .CP(clk), 
        .Q(\stage_2_retimer[5][8] ) );
  DFQD1 \stage_2_retimer_reg[5][7]  ( .D(\stage_2_output[5][7] ), .CP(clk), 
        .Q(\stage_2_retimer[5][7] ) );
  DFQD1 \stage_2_retimer_reg[5][6]  ( .D(\stage_2_output[5][6] ), .CP(clk), 
        .Q(\stage_2_retimer[5][6] ) );
  DFQD1 \stage_2_retimer_reg[5][5]  ( .D(\stage_2_output[5][5] ), .CP(clk), 
        .Q(\stage_2_retimer[5][5] ) );
  DFQD1 \stage_2_retimer_reg[5][4]  ( .D(\stage_2_output[5][4] ), .CP(clk), 
        .Q(\stage_2_retimer[5][4] ) );
  DFQD1 \stage_2_retimer_reg[5][3]  ( .D(\stage_2_output[5][3] ), .CP(clk), 
        .Q(\stage_2_retimer[5][3] ) );
  DFQD1 \stage_2_retimer_reg[5][2]  ( .D(\stage_2_output[5][2] ), .CP(clk), 
        .Q(\stage_2_retimer[5][2] ) );
  DFQD1 \stage_2_retimer_reg[5][1]  ( .D(\stage_2_output[5][1] ), .CP(clk), 
        .Q(\stage_2_retimer[5][1] ) );
  DFQD1 \stage_2_retimer_reg[5][0]  ( .D(\stage_2_output[5][0] ), .CP(clk), 
        .Q(\stage_2_retimer[5][0] ) );
  DFQD1 \stage_2_retimer_reg[4][19]  ( .D(\stage_2_output[4][19] ), .CP(clk), 
        .Q(\stage_2_retimer[4][19] ) );
  DFQD1 \stage_2_retimer_reg[4][18]  ( .D(\stage_2_output[4][18] ), .CP(clk), 
        .Q(\stage_2_retimer[4][18] ) );
  DFQD1 \stage_2_retimer_reg[4][17]  ( .D(\stage_2_output[4][17] ), .CP(clk), 
        .Q(\stage_2_retimer[4][17] ) );
  DFQD1 \stage_2_retimer_reg[4][16]  ( .D(\stage_2_output[4][16] ), .CP(clk), 
        .Q(\stage_2_retimer[4][16] ) );
  DFQD1 \stage_2_retimer_reg[4][15]  ( .D(\stage_2_output[4][15] ), .CP(clk), 
        .Q(\stage_2_retimer[4][15] ) );
  DFQD1 \stage_2_retimer_reg[4][14]  ( .D(\stage_2_output[4][14] ), .CP(clk), 
        .Q(\stage_2_retimer[4][14] ) );
  DFQD1 \stage_2_retimer_reg[4][13]  ( .D(\stage_2_output[4][13] ), .CP(clk), 
        .Q(\stage_2_retimer[4][13] ) );
  DFQD1 \stage_2_retimer_reg[4][12]  ( .D(\stage_2_output[4][12] ), .CP(clk), 
        .Q(\stage_2_retimer[4][12] ) );
  DFQD1 \stage_2_retimer_reg[4][11]  ( .D(\stage_2_output[4][11] ), .CP(clk), 
        .Q(\stage_2_retimer[4][11] ) );
  DFQD1 \stage_2_retimer_reg[4][10]  ( .D(\stage_2_output[4][10] ), .CP(clk), 
        .Q(\stage_2_retimer[4][10] ) );
  DFQD1 \stage_2_retimer_reg[4][9]  ( .D(\stage_2_output[4][9] ), .CP(clk), 
        .Q(\stage_2_retimer[4][9] ) );
  DFQD1 \stage_2_retimer_reg[4][8]  ( .D(\stage_2_output[4][8] ), .CP(clk), 
        .Q(\stage_2_retimer[4][8] ) );
  DFQD1 \stage_2_retimer_reg[4][7]  ( .D(\stage_2_output[4][7] ), .CP(clk), 
        .Q(\stage_2_retimer[4][7] ) );
  DFQD1 \stage_2_retimer_reg[4][6]  ( .D(\stage_2_output[4][6] ), .CP(clk), 
        .Q(\stage_2_retimer[4][6] ) );
  DFQD1 \stage_2_retimer_reg[4][5]  ( .D(\stage_2_output[4][5] ), .CP(clk), 
        .Q(\stage_2_retimer[4][5] ) );
  DFQD1 \stage_2_retimer_reg[4][4]  ( .D(\stage_2_output[4][4] ), .CP(clk), 
        .Q(\stage_2_retimer[4][4] ) );
  DFQD1 \stage_2_retimer_reg[4][3]  ( .D(\stage_2_output[4][3] ), .CP(clk), 
        .Q(\stage_2_retimer[4][3] ) );
  DFQD1 \stage_2_retimer_reg[4][2]  ( .D(\stage_2_output[4][2] ), .CP(clk), 
        .Q(\stage_2_retimer[4][2] ) );
  DFQD1 \stage_2_retimer_reg[4][1]  ( .D(\stage_2_output[4][1] ), .CP(clk), 
        .Q(\stage_2_retimer[4][1] ) );
  DFQD1 \stage_2_retimer_reg[4][0]  ( .D(\stage_2_output[4][0] ), .CP(clk), 
        .Q(\stage_2_retimer[4][0] ) );
  DFQD1 \stage_2_retimer_reg[3][19]  ( .D(\stage_2_output[3][19] ), .CP(clk), 
        .Q(\stage_2_retimer[3][19] ) );
  DFQD1 \stage_2_retimer_reg[3][18]  ( .D(\stage_2_output[3][18] ), .CP(clk), 
        .Q(\stage_2_retimer[3][18] ) );
  DFQD1 \stage_2_retimer_reg[3][17]  ( .D(\stage_2_output[3][17] ), .CP(clk), 
        .Q(\stage_2_retimer[3][17] ) );
  DFQD1 \stage_2_retimer_reg[3][16]  ( .D(\stage_2_output[3][16] ), .CP(clk), 
        .Q(\stage_2_retimer[3][16] ) );
  DFQD1 \stage_2_retimer_reg[3][15]  ( .D(\stage_2_output[3][15] ), .CP(clk), 
        .Q(\stage_2_retimer[3][15] ) );
  DFQD1 \stage_2_retimer_reg[3][14]  ( .D(\stage_2_output[3][14] ), .CP(clk), 
        .Q(\stage_2_retimer[3][14] ) );
  DFQD1 \stage_2_retimer_reg[3][13]  ( .D(\stage_2_output[3][13] ), .CP(clk), 
        .Q(\stage_2_retimer[3][13] ) );
  DFQD1 \stage_2_retimer_reg[3][12]  ( .D(\stage_2_output[3][12] ), .CP(clk), 
        .Q(\stage_2_retimer[3][12] ) );
  DFQD1 \stage_2_retimer_reg[3][11]  ( .D(\stage_2_output[3][11] ), .CP(clk), 
        .Q(\stage_2_retimer[3][11] ) );
  DFQD1 \stage_2_retimer_reg[3][10]  ( .D(\stage_2_output[3][10] ), .CP(clk), 
        .Q(\stage_2_retimer[3][10] ) );
  DFQD1 \stage_2_retimer_reg[3][9]  ( .D(\stage_2_output[3][9] ), .CP(clk), 
        .Q(\stage_2_retimer[3][9] ) );
  DFQD1 \stage_2_retimer_reg[3][8]  ( .D(\stage_2_output[3][8] ), .CP(clk), 
        .Q(\stage_2_retimer[3][8] ) );
  DFQD1 \stage_2_retimer_reg[3][7]  ( .D(\stage_2_output[3][7] ), .CP(clk), 
        .Q(\stage_2_retimer[3][7] ) );
  DFQD1 \stage_2_retimer_reg[3][6]  ( .D(\stage_2_output[3][6] ), .CP(clk), 
        .Q(\stage_2_retimer[3][6] ) );
  DFQD1 \stage_2_retimer_reg[3][5]  ( .D(\stage_2_output[3][5] ), .CP(clk), 
        .Q(\stage_2_retimer[3][5] ) );
  DFQD1 \stage_2_retimer_reg[3][4]  ( .D(\stage_2_output[3][4] ), .CP(clk), 
        .Q(\stage_2_retimer[3][4] ) );
  DFQD1 \stage_2_retimer_reg[3][3]  ( .D(\stage_2_output[3][3] ), .CP(clk), 
        .Q(\stage_2_retimer[3][3] ) );
  DFQD1 \stage_2_retimer_reg[3][2]  ( .D(\stage_2_output[3][2] ), .CP(clk), 
        .Q(\stage_2_retimer[3][2] ) );
  DFQD1 \stage_2_retimer_reg[3][1]  ( .D(\stage_2_output[3][1] ), .CP(clk), 
        .Q(\stage_2_retimer[3][1] ) );
  DFQD1 \stage_2_retimer_reg[3][0]  ( .D(\stage_2_output[3][0] ), .CP(clk), 
        .Q(\stage_2_retimer[3][0] ) );
  DFQD1 \stage_2_retimer_reg[2][19]  ( .D(\stage_2_output[2][19] ), .CP(clk), 
        .Q(\stage_2_retimer[2][19] ) );
  DFQD1 \stage_2_retimer_reg[2][18]  ( .D(\stage_2_output[2][18] ), .CP(clk), 
        .Q(\stage_2_retimer[2][18] ) );
  DFQD1 \stage_2_retimer_reg[2][17]  ( .D(\stage_2_output[2][17] ), .CP(clk), 
        .Q(\stage_2_retimer[2][17] ) );
  DFQD1 \stage_2_retimer_reg[2][16]  ( .D(\stage_2_output[2][16] ), .CP(clk), 
        .Q(\stage_2_retimer[2][16] ) );
  DFQD1 \stage_2_retimer_reg[2][15]  ( .D(\stage_2_output[2][15] ), .CP(clk), 
        .Q(\stage_2_retimer[2][15] ) );
  DFQD1 \stage_2_retimer_reg[2][14]  ( .D(\stage_2_output[2][14] ), .CP(clk), 
        .Q(\stage_2_retimer[2][14] ) );
  DFQD1 \stage_2_retimer_reg[2][13]  ( .D(\stage_2_output[2][13] ), .CP(clk), 
        .Q(\stage_2_retimer[2][13] ) );
  DFQD1 \stage_2_retimer_reg[2][12]  ( .D(\stage_2_output[2][12] ), .CP(clk), 
        .Q(\stage_2_retimer[2][12] ) );
  DFQD1 \stage_2_retimer_reg[2][11]  ( .D(\stage_2_output[2][11] ), .CP(clk), 
        .Q(\stage_2_retimer[2][11] ) );
  DFQD1 \stage_2_retimer_reg[2][10]  ( .D(\stage_2_output[2][10] ), .CP(clk), 
        .Q(\stage_2_retimer[2][10] ) );
  DFQD1 \stage_2_retimer_reg[2][9]  ( .D(\stage_2_output[2][9] ), .CP(clk), 
        .Q(\stage_2_retimer[2][9] ) );
  DFQD1 \stage_2_retimer_reg[2][8]  ( .D(\stage_2_output[2][8] ), .CP(clk), 
        .Q(\stage_2_retimer[2][8] ) );
  DFQD1 \stage_2_retimer_reg[2][7]  ( .D(\stage_2_output[2][7] ), .CP(clk), 
        .Q(\stage_2_retimer[2][7] ) );
  DFQD1 \stage_2_retimer_reg[2][6]  ( .D(\stage_2_output[2][6] ), .CP(clk), 
        .Q(\stage_2_retimer[2][6] ) );
  DFQD1 \stage_2_retimer_reg[2][5]  ( .D(\stage_2_output[2][5] ), .CP(clk), 
        .Q(\stage_2_retimer[2][5] ) );
  DFQD1 \stage_2_retimer_reg[2][4]  ( .D(\stage_2_output[2][4] ), .CP(clk), 
        .Q(\stage_2_retimer[2][4] ) );
  DFQD1 \stage_2_retimer_reg[2][3]  ( .D(\stage_2_output[2][3] ), .CP(clk), 
        .Q(\stage_2_retimer[2][3] ) );
  DFQD1 \stage_2_retimer_reg[2][2]  ( .D(\stage_2_output[2][2] ), .CP(clk), 
        .Q(\stage_2_retimer[2][2] ) );
  DFQD1 \stage_2_retimer_reg[2][1]  ( .D(\stage_2_output[2][1] ), .CP(clk), 
        .Q(\stage_2_retimer[2][1] ) );
  DFQD1 \stage_2_retimer_reg[2][0]  ( .D(\stage_2_output[2][0] ), .CP(clk), 
        .Q(\stage_2_retimer[2][0] ) );
  DFQD1 \stage_2_retimer_reg[1][19]  ( .D(\stage_2_output[1][19] ), .CP(clk), 
        .Q(\stage_2_retimer[1][19] ) );
  DFQD1 \stage_2_retimer_reg[1][18]  ( .D(\stage_2_output[1][18] ), .CP(clk), 
        .Q(\stage_2_retimer[1][18] ) );
  DFQD1 \stage_2_retimer_reg[1][17]  ( .D(\stage_2_output[1][17] ), .CP(clk), 
        .Q(\stage_2_retimer[1][17] ) );
  DFQD1 \stage_2_retimer_reg[1][16]  ( .D(\stage_2_output[1][16] ), .CP(clk), 
        .Q(\stage_2_retimer[1][16] ) );
  DFQD1 \stage_2_retimer_reg[1][15]  ( .D(\stage_2_output[1][15] ), .CP(clk), 
        .Q(\stage_2_retimer[1][15] ) );
  DFQD1 \stage_2_retimer_reg[1][14]  ( .D(\stage_2_output[1][14] ), .CP(clk), 
        .Q(\stage_2_retimer[1][14] ) );
  DFQD1 \stage_2_retimer_reg[1][13]  ( .D(\stage_2_output[1][13] ), .CP(clk), 
        .Q(\stage_2_retimer[1][13] ) );
  DFQD1 \stage_2_retimer_reg[1][12]  ( .D(\stage_2_output[1][12] ), .CP(clk), 
        .Q(\stage_2_retimer[1][12] ) );
  DFQD1 \stage_2_retimer_reg[1][11]  ( .D(\stage_2_output[1][11] ), .CP(clk), 
        .Q(\stage_2_retimer[1][11] ) );
  DFQD1 \stage_2_retimer_reg[1][10]  ( .D(\stage_2_output[1][10] ), .CP(clk), 
        .Q(\stage_2_retimer[1][10] ) );
  DFQD1 \stage_2_retimer_reg[1][9]  ( .D(\stage_2_output[1][9] ), .CP(clk), 
        .Q(\stage_2_retimer[1][9] ) );
  DFQD1 \stage_2_retimer_reg[1][8]  ( .D(\stage_2_output[1][8] ), .CP(clk), 
        .Q(\stage_2_retimer[1][8] ) );
  DFQD1 \stage_2_retimer_reg[1][7]  ( .D(\stage_2_output[1][7] ), .CP(clk), 
        .Q(\stage_2_retimer[1][7] ) );
  DFQD1 \stage_2_retimer_reg[1][6]  ( .D(\stage_2_output[1][6] ), .CP(clk), 
        .Q(\stage_2_retimer[1][6] ) );
  DFQD1 \stage_2_retimer_reg[1][5]  ( .D(\stage_2_output[1][5] ), .CP(clk), 
        .Q(\stage_2_retimer[1][5] ) );
  DFQD1 \stage_2_retimer_reg[1][4]  ( .D(\stage_2_output[1][4] ), .CP(clk), 
        .Q(\stage_2_retimer[1][4] ) );
  DFQD1 \stage_2_retimer_reg[1][3]  ( .D(\stage_2_output[1][3] ), .CP(clk), 
        .Q(\stage_2_retimer[1][3] ) );
  DFQD1 \stage_2_retimer_reg[1][2]  ( .D(\stage_2_output[1][2] ), .CP(clk), 
        .Q(\stage_2_retimer[1][2] ) );
  DFQD1 \stage_2_retimer_reg[1][1]  ( .D(\stage_2_output[1][1] ), .CP(clk), 
        .Q(\stage_2_retimer[1][1] ) );
  DFQD1 \stage_2_retimer_reg[1][0]  ( .D(\stage_2_output[1][0] ), .CP(clk), 
        .Q(\stage_2_retimer[1][0] ) );
  DFQD1 \stage_2_retimer_reg[0][19]  ( .D(\stage_2_output[0][19] ), .CP(clk), 
        .Q(\stage_2_retimer[0][19] ) );
  DFQD1 \stage_2_retimer_reg[0][18]  ( .D(\stage_2_output[0][18] ), .CP(clk), 
        .Q(\stage_2_retimer[0][18] ) );
  DFQD1 \stage_2_retimer_reg[0][17]  ( .D(\stage_2_output[0][17] ), .CP(clk), 
        .Q(\stage_2_retimer[0][17] ) );
  DFQD1 \stage_2_retimer_reg[0][16]  ( .D(\stage_2_output[0][16] ), .CP(clk), 
        .Q(\stage_2_retimer[0][16] ) );
  DFQD1 \stage_2_retimer_reg[0][15]  ( .D(\stage_2_output[0][15] ), .CP(clk), 
        .Q(\stage_2_retimer[0][15] ) );
  DFQD1 \stage_2_retimer_reg[0][14]  ( .D(\stage_2_output[0][14] ), .CP(clk), 
        .Q(\stage_2_retimer[0][14] ) );
  DFQD1 \stage_2_retimer_reg[0][13]  ( .D(\stage_2_output[0][13] ), .CP(clk), 
        .Q(\stage_2_retimer[0][13] ) );
  DFQD1 \stage_2_retimer_reg[0][12]  ( .D(\stage_2_output[0][12] ), .CP(clk), 
        .Q(\stage_2_retimer[0][12] ) );
  DFQD1 \stage_2_retimer_reg[0][11]  ( .D(\stage_2_output[0][11] ), .CP(clk), 
        .Q(\stage_2_retimer[0][11] ) );
  DFQD1 \stage_2_retimer_reg[0][10]  ( .D(\stage_2_output[0][10] ), .CP(clk), 
        .Q(\stage_2_retimer[0][10] ) );
  DFQD1 \stage_2_retimer_reg[0][9]  ( .D(\stage_2_output[0][9] ), .CP(clk), 
        .Q(\stage_2_retimer[0][9] ) );
  DFQD1 \stage_2_retimer_reg[0][8]  ( .D(\stage_2_output[0][8] ), .CP(clk), 
        .Q(\stage_2_retimer[0][8] ) );
  DFQD1 \stage_2_retimer_reg[0][7]  ( .D(\stage_2_output[0][7] ), .CP(clk), 
        .Q(\stage_2_retimer[0][7] ) );
  DFQD1 \stage_2_retimer_reg[0][6]  ( .D(\stage_2_output[0][6] ), .CP(clk), 
        .Q(\stage_2_retimer[0][6] ) );
  DFQD1 \stage_2_retimer_reg[0][5]  ( .D(\stage_2_output[0][5] ), .CP(clk), 
        .Q(\stage_2_retimer[0][5] ) );
  DFQD1 \stage_2_retimer_reg[0][4]  ( .D(\stage_2_output[0][4] ), .CP(clk), 
        .Q(\stage_2_retimer[0][4] ) );
  DFQD1 \stage_2_retimer_reg[0][3]  ( .D(\stage_2_output[0][3] ), .CP(clk), 
        .Q(\stage_2_retimer[0][3] ) );
  DFQD1 \stage_2_retimer_reg[0][2]  ( .D(\stage_2_output[0][2] ), .CP(clk), 
        .Q(\stage_2_retimer[0][2] ) );
  DFQD1 \stage_2_retimer_reg[0][1]  ( .D(\stage_2_output[0][1] ), .CP(clk), 
        .Q(\stage_2_retimer[0][1] ) );
  DFQD1 \stage_2_retimer_reg[0][0]  ( .D(\stage_2_output[0][0] ), .CP(clk), 
        .Q(\stage_2_retimer[0][0] ) );
  DFQD1 \stage_3_retimer_reg[7][19]  ( .D(\stage_3_output[7][19] ), .CP(clk), 
        .Q(\stage_3_retimer[7][19] ) );
  DFQD1 \stage_3_retimer_reg[7][18]  ( .D(\stage_3_output[7][18] ), .CP(clk), 
        .Q(\stage_3_retimer[7][18] ) );
  DFQD1 \stage_3_retimer_reg[7][17]  ( .D(\stage_3_output[7][17] ), .CP(clk), 
        .Q(\stage_3_retimer[7][17] ) );
  DFQD1 \stage_3_retimer_reg[7][16]  ( .D(\stage_3_output[7][16] ), .CP(clk), 
        .Q(\stage_3_retimer[7][16] ) );
  DFQD1 \stage_3_retimer_reg[7][15]  ( .D(\stage_3_output[7][15] ), .CP(clk), 
        .Q(\stage_3_retimer[7][15] ) );
  DFQD1 \stage_3_retimer_reg[7][14]  ( .D(\stage_3_output[7][14] ), .CP(clk), 
        .Q(\stage_3_retimer[7][14] ) );
  DFQD1 \stage_3_retimer_reg[7][13]  ( .D(\stage_3_output[7][13] ), .CP(clk), 
        .Q(\stage_3_retimer[7][13] ) );
  DFQD1 \stage_3_retimer_reg[7][12]  ( .D(\stage_3_output[7][12] ), .CP(clk), 
        .Q(\stage_3_retimer[7][12] ) );
  DFQD1 \stage_3_retimer_reg[7][11]  ( .D(\stage_3_output[7][11] ), .CP(clk), 
        .Q(\stage_3_retimer[7][11] ) );
  DFQD1 \stage_3_retimer_reg[7][10]  ( .D(\stage_3_output[7][10] ), .CP(clk), 
        .Q(\stage_3_retimer[7][10] ) );
  DFQD1 \stage_3_retimer_reg[7][9]  ( .D(\stage_3_output[7][9] ), .CP(clk), 
        .Q(\stage_3_retimer[7][9] ) );
  DFQD1 \stage_3_retimer_reg[7][8]  ( .D(\stage_3_output[7][8] ), .CP(clk), 
        .Q(\stage_3_retimer[7][8] ) );
  DFQD1 \stage_3_retimer_reg[7][7]  ( .D(\stage_3_output[7][7] ), .CP(clk), 
        .Q(\stage_3_retimer[7][7] ) );
  DFQD1 \stage_3_retimer_reg[7][6]  ( .D(\stage_3_output[7][6] ), .CP(clk), 
        .Q(\stage_3_retimer[7][6] ) );
  DFQD1 \stage_3_retimer_reg[7][5]  ( .D(\stage_3_output[7][5] ), .CP(clk), 
        .Q(\stage_3_retimer[7][5] ) );
  DFQD1 \stage_3_retimer_reg[7][4]  ( .D(\stage_3_output[7][4] ), .CP(clk), 
        .Q(\stage_3_retimer[7][4] ) );
  DFQD1 \stage_3_retimer_reg[7][3]  ( .D(\stage_3_output[7][3] ), .CP(clk), 
        .Q(\stage_3_retimer[7][3] ) );
  DFQD1 \stage_3_retimer_reg[7][2]  ( .D(\stage_3_output[7][2] ), .CP(clk), 
        .Q(\stage_3_retimer[7][2] ) );
  DFQD1 \stage_3_retimer_reg[7][1]  ( .D(\stage_3_output[7][1] ), .CP(clk), 
        .Q(\stage_3_retimer[7][1] ) );
  DFQD1 \stage_3_retimer_reg[7][0]  ( .D(\stage_3_output[7][0] ), .CP(clk), 
        .Q(\stage_3_retimer[7][0] ) );
  DFQD1 \stage_3_retimer_reg[6][19]  ( .D(\stage_3_output[6][19] ), .CP(clk), 
        .Q(\stage_3_retimer[6][19] ) );
  DFQD1 \stage_3_retimer_reg[6][18]  ( .D(\stage_3_output[6][18] ), .CP(clk), 
        .Q(\stage_3_retimer[6][18] ) );
  DFQD1 \stage_3_retimer_reg[6][17]  ( .D(\stage_3_output[6][17] ), .CP(clk), 
        .Q(\stage_3_retimer[6][17] ) );
  DFQD1 \stage_3_retimer_reg[6][16]  ( .D(\stage_3_output[6][16] ), .CP(clk), 
        .Q(\stage_3_retimer[6][16] ) );
  DFQD1 \stage_3_retimer_reg[6][15]  ( .D(\stage_3_output[6][15] ), .CP(clk), 
        .Q(\stage_3_retimer[6][15] ) );
  DFQD1 \stage_3_retimer_reg[6][14]  ( .D(\stage_3_output[6][14] ), .CP(clk), 
        .Q(\stage_3_retimer[6][14] ) );
  DFQD1 \stage_3_retimer_reg[6][13]  ( .D(\stage_3_output[6][13] ), .CP(clk), 
        .Q(\stage_3_retimer[6][13] ) );
  DFQD1 \stage_3_retimer_reg[6][12]  ( .D(\stage_3_output[6][12] ), .CP(clk), 
        .Q(\stage_3_retimer[6][12] ) );
  DFQD1 \stage_3_retimer_reg[6][11]  ( .D(\stage_3_output[6][11] ), .CP(clk), 
        .Q(\stage_3_retimer[6][11] ) );
  DFQD1 \stage_3_retimer_reg[6][10]  ( .D(\stage_3_output[6][10] ), .CP(clk), 
        .Q(\stage_3_retimer[6][10] ) );
  DFQD1 \stage_3_retimer_reg[6][9]  ( .D(\stage_3_output[6][9] ), .CP(clk), 
        .Q(\stage_3_retimer[6][9] ) );
  DFQD1 \stage_3_retimer_reg[6][8]  ( .D(\stage_3_output[6][8] ), .CP(clk), 
        .Q(\stage_3_retimer[6][8] ) );
  DFQD1 \stage_3_retimer_reg[6][7]  ( .D(\stage_3_output[6][7] ), .CP(clk), 
        .Q(\stage_3_retimer[6][7] ) );
  DFQD1 \stage_3_retimer_reg[6][6]  ( .D(\stage_3_output[6][6] ), .CP(clk), 
        .Q(\stage_3_retimer[6][6] ) );
  DFQD1 \stage_3_retimer_reg[6][5]  ( .D(\stage_3_output[6][5] ), .CP(clk), 
        .Q(\stage_3_retimer[6][5] ) );
  DFQD1 \stage_3_retimer_reg[6][4]  ( .D(\stage_3_output[6][4] ), .CP(clk), 
        .Q(\stage_3_retimer[6][4] ) );
  DFQD1 \stage_3_retimer_reg[6][3]  ( .D(\stage_3_output[6][3] ), .CP(clk), 
        .Q(\stage_3_retimer[6][3] ) );
  DFQD1 \stage_3_retimer_reg[6][2]  ( .D(\stage_3_output[6][2] ), .CP(clk), 
        .Q(\stage_3_retimer[6][2] ) );
  DFQD1 \stage_3_retimer_reg[6][1]  ( .D(\stage_3_output[6][1] ), .CP(clk), 
        .Q(\stage_3_retimer[6][1] ) );
  DFQD1 \stage_3_retimer_reg[6][0]  ( .D(\stage_3_output[6][0] ), .CP(clk), 
        .Q(\stage_3_retimer[6][0] ) );
  DFQD1 \stage_3_retimer_reg[5][19]  ( .D(\stage_3_output[5][19] ), .CP(clk), 
        .Q(\stage_3_retimer[5][19] ) );
  DFQD1 \stage_3_retimer_reg[5][18]  ( .D(\stage_3_output[5][18] ), .CP(clk), 
        .Q(\stage_3_retimer[5][18] ) );
  DFQD1 \stage_3_retimer_reg[5][17]  ( .D(\stage_3_output[5][17] ), .CP(clk), 
        .Q(\stage_3_retimer[5][17] ) );
  DFQD1 \stage_3_retimer_reg[5][16]  ( .D(\stage_3_output[5][16] ), .CP(clk), 
        .Q(\stage_3_retimer[5][16] ) );
  DFQD1 \stage_3_retimer_reg[5][15]  ( .D(\stage_3_output[5][15] ), .CP(clk), 
        .Q(\stage_3_retimer[5][15] ) );
  DFQD1 \stage_3_retimer_reg[5][14]  ( .D(\stage_3_output[5][14] ), .CP(clk), 
        .Q(\stage_3_retimer[5][14] ) );
  DFQD1 \stage_3_retimer_reg[5][13]  ( .D(\stage_3_output[5][13] ), .CP(clk), 
        .Q(\stage_3_retimer[5][13] ) );
  DFQD1 \stage_3_retimer_reg[5][12]  ( .D(\stage_3_output[5][12] ), .CP(clk), 
        .Q(\stage_3_retimer[5][12] ) );
  DFQD1 \stage_3_retimer_reg[5][11]  ( .D(\stage_3_output[5][11] ), .CP(clk), 
        .Q(\stage_3_retimer[5][11] ) );
  DFQD1 \stage_3_retimer_reg[5][10]  ( .D(\stage_3_output[5][10] ), .CP(clk), 
        .Q(\stage_3_retimer[5][10] ) );
  DFQD1 \stage_3_retimer_reg[5][9]  ( .D(\stage_3_output[5][9] ), .CP(clk), 
        .Q(\stage_3_retimer[5][9] ) );
  DFQD1 \stage_3_retimer_reg[5][8]  ( .D(\stage_3_output[5][8] ), .CP(clk), 
        .Q(\stage_3_retimer[5][8] ) );
  DFQD1 \stage_3_retimer_reg[5][7]  ( .D(\stage_3_output[5][7] ), .CP(clk), 
        .Q(\stage_3_retimer[5][7] ) );
  DFQD1 \stage_3_retimer_reg[5][6]  ( .D(\stage_3_output[5][6] ), .CP(clk), 
        .Q(\stage_3_retimer[5][6] ) );
  DFQD1 \stage_3_retimer_reg[5][5]  ( .D(\stage_3_output[5][5] ), .CP(clk), 
        .Q(\stage_3_retimer[5][5] ) );
  DFQD1 \stage_3_retimer_reg[5][4]  ( .D(\stage_3_output[5][4] ), .CP(clk), 
        .Q(\stage_3_retimer[5][4] ) );
  DFQD1 \stage_3_retimer_reg[5][3]  ( .D(\stage_3_output[5][3] ), .CP(clk), 
        .Q(\stage_3_retimer[5][3] ) );
  DFQD1 \stage_3_retimer_reg[5][2]  ( .D(\stage_3_output[5][2] ), .CP(clk), 
        .Q(\stage_3_retimer[5][2] ) );
  DFQD1 \stage_3_retimer_reg[5][1]  ( .D(\stage_3_output[5][1] ), .CP(clk), 
        .Q(\stage_3_retimer[5][1] ) );
  DFQD1 \stage_3_retimer_reg[5][0]  ( .D(\stage_3_output[5][0] ), .CP(clk), 
        .Q(\stage_3_retimer[5][0] ) );
  DFQD1 \stage_3_retimer_reg[4][19]  ( .D(\stage_3_output[4][19] ), .CP(clk), 
        .Q(\stage_3_retimer[4][19] ) );
  DFQD1 \stage_3_retimer_reg[4][18]  ( .D(\stage_3_output[4][18] ), .CP(clk), 
        .Q(\stage_3_retimer[4][18] ) );
  DFQD1 \stage_3_retimer_reg[4][17]  ( .D(\stage_3_output[4][17] ), .CP(clk), 
        .Q(\stage_3_retimer[4][17] ) );
  DFQD1 \stage_3_retimer_reg[4][16]  ( .D(\stage_3_output[4][16] ), .CP(clk), 
        .Q(\stage_3_retimer[4][16] ) );
  DFQD1 \stage_3_retimer_reg[4][15]  ( .D(\stage_3_output[4][15] ), .CP(clk), 
        .Q(\stage_3_retimer[4][15] ) );
  DFQD1 \stage_3_retimer_reg[4][14]  ( .D(\stage_3_output[4][14] ), .CP(clk), 
        .Q(\stage_3_retimer[4][14] ) );
  DFQD1 \stage_3_retimer_reg[4][13]  ( .D(\stage_3_output[4][13] ), .CP(clk), 
        .Q(\stage_3_retimer[4][13] ) );
  DFQD1 \stage_3_retimer_reg[4][12]  ( .D(\stage_3_output[4][12] ), .CP(clk), 
        .Q(\stage_3_retimer[4][12] ) );
  DFQD1 \stage_3_retimer_reg[4][11]  ( .D(\stage_3_output[4][11] ), .CP(clk), 
        .Q(\stage_3_retimer[4][11] ) );
  DFQD1 \stage_3_retimer_reg[4][10]  ( .D(\stage_3_output[4][10] ), .CP(clk), 
        .Q(\stage_3_retimer[4][10] ) );
  DFQD1 \stage_3_retimer_reg[4][9]  ( .D(\stage_3_output[4][9] ), .CP(clk), 
        .Q(\stage_3_retimer[4][9] ) );
  DFQD1 \stage_3_retimer_reg[4][8]  ( .D(\stage_3_output[4][8] ), .CP(clk), 
        .Q(\stage_3_retimer[4][8] ) );
  DFQD1 \stage_3_retimer_reg[4][7]  ( .D(\stage_3_output[4][7] ), .CP(clk), 
        .Q(\stage_3_retimer[4][7] ) );
  DFQD1 \stage_3_retimer_reg[4][6]  ( .D(\stage_3_output[4][6] ), .CP(clk), 
        .Q(\stage_3_retimer[4][6] ) );
  DFQD1 \stage_3_retimer_reg[4][5]  ( .D(\stage_3_output[4][5] ), .CP(clk), 
        .Q(\stage_3_retimer[4][5] ) );
  DFQD1 \stage_3_retimer_reg[4][4]  ( .D(\stage_3_output[4][4] ), .CP(clk), 
        .Q(\stage_3_retimer[4][4] ) );
  DFQD1 \stage_3_retimer_reg[4][3]  ( .D(\stage_3_output[4][3] ), .CP(clk), 
        .Q(\stage_3_retimer[4][3] ) );
  DFQD1 \stage_3_retimer_reg[4][2]  ( .D(\stage_3_output[4][2] ), .CP(clk), 
        .Q(\stage_3_retimer[4][2] ) );
  DFQD1 \stage_3_retimer_reg[4][1]  ( .D(\stage_3_output[4][1] ), .CP(clk), 
        .Q(\stage_3_retimer[4][1] ) );
  DFQD1 \stage_3_retimer_reg[4][0]  ( .D(\stage_3_output[4][0] ), .CP(clk), 
        .Q(\stage_3_retimer[4][0] ) );
  DFQD1 \stage_3_retimer_reg[3][19]  ( .D(\stage_3_output[3][19] ), .CP(clk), 
        .Q(\stage_3_retimer[3][19] ) );
  DFQD1 \stage_3_retimer_reg[3][18]  ( .D(\stage_3_output[3][18] ), .CP(clk), 
        .Q(\stage_3_retimer[3][18] ) );
  DFQD1 \stage_3_retimer_reg[3][17]  ( .D(\stage_3_output[3][17] ), .CP(clk), 
        .Q(\stage_3_retimer[3][17] ) );
  DFQD1 \stage_3_retimer_reg[3][16]  ( .D(\stage_3_output[3][16] ), .CP(clk), 
        .Q(\stage_3_retimer[3][16] ) );
  DFQD1 \stage_3_retimer_reg[3][15]  ( .D(\stage_3_output[3][15] ), .CP(clk), 
        .Q(\stage_3_retimer[3][15] ) );
  DFQD1 \stage_3_retimer_reg[3][14]  ( .D(\stage_3_output[3][14] ), .CP(clk), 
        .Q(\stage_3_retimer[3][14] ) );
  DFQD1 \stage_3_retimer_reg[3][13]  ( .D(\stage_3_output[3][13] ), .CP(clk), 
        .Q(\stage_3_retimer[3][13] ) );
  DFQD1 \stage_3_retimer_reg[3][12]  ( .D(\stage_3_output[3][12] ), .CP(clk), 
        .Q(\stage_3_retimer[3][12] ) );
  DFQD1 \stage_3_retimer_reg[3][11]  ( .D(\stage_3_output[3][11] ), .CP(clk), 
        .Q(\stage_3_retimer[3][11] ) );
  DFQD1 \stage_3_retimer_reg[3][10]  ( .D(\stage_3_output[3][10] ), .CP(clk), 
        .Q(\stage_3_retimer[3][10] ) );
  DFQD1 \stage_3_retimer_reg[3][9]  ( .D(\stage_3_output[3][9] ), .CP(clk), 
        .Q(\stage_3_retimer[3][9] ) );
  DFQD1 \stage_3_retimer_reg[3][8]  ( .D(\stage_3_output[3][8] ), .CP(clk), 
        .Q(\stage_3_retimer[3][8] ) );
  DFQD1 \stage_3_retimer_reg[3][7]  ( .D(\stage_3_output[3][7] ), .CP(clk), 
        .Q(\stage_3_retimer[3][7] ) );
  DFQD1 \stage_3_retimer_reg[3][6]  ( .D(\stage_3_output[3][6] ), .CP(clk), 
        .Q(\stage_3_retimer[3][6] ) );
  DFQD1 \stage_3_retimer_reg[3][5]  ( .D(\stage_3_output[3][5] ), .CP(clk), 
        .Q(\stage_3_retimer[3][5] ) );
  DFQD1 \stage_3_retimer_reg[3][4]  ( .D(\stage_3_output[3][4] ), .CP(clk), 
        .Q(\stage_3_retimer[3][4] ) );
  DFQD1 \stage_3_retimer_reg[3][3]  ( .D(\stage_3_output[3][3] ), .CP(clk), 
        .Q(\stage_3_retimer[3][3] ) );
  DFQD1 \stage_3_retimer_reg[3][2]  ( .D(\stage_3_output[3][2] ), .CP(clk), 
        .Q(\stage_3_retimer[3][2] ) );
  DFQD1 \stage_3_retimer_reg[3][1]  ( .D(\stage_3_output[3][1] ), .CP(clk), 
        .Q(\stage_3_retimer[3][1] ) );
  DFQD1 \stage_3_retimer_reg[3][0]  ( .D(\stage_3_output[3][0] ), .CP(clk), 
        .Q(\stage_3_retimer[3][0] ) );
  DFQD1 \stage_3_retimer_reg[2][19]  ( .D(\stage_3_output[2][19] ), .CP(clk), 
        .Q(\stage_3_retimer[2][19] ) );
  DFQD1 \stage_3_retimer_reg[2][18]  ( .D(\stage_3_output[2][18] ), .CP(clk), 
        .Q(\stage_3_retimer[2][18] ) );
  DFQD1 \stage_3_retimer_reg[2][17]  ( .D(\stage_3_output[2][17] ), .CP(clk), 
        .Q(\stage_3_retimer[2][17] ) );
  DFQD1 \stage_3_retimer_reg[2][16]  ( .D(\stage_3_output[2][16] ), .CP(clk), 
        .Q(\stage_3_retimer[2][16] ) );
  DFQD1 \stage_3_retimer_reg[2][15]  ( .D(\stage_3_output[2][15] ), .CP(clk), 
        .Q(\stage_3_retimer[2][15] ) );
  DFQD1 \stage_3_retimer_reg[2][14]  ( .D(\stage_3_output[2][14] ), .CP(clk), 
        .Q(\stage_3_retimer[2][14] ) );
  DFQD1 \stage_3_retimer_reg[2][13]  ( .D(\stage_3_output[2][13] ), .CP(clk), 
        .Q(\stage_3_retimer[2][13] ) );
  DFQD1 \stage_3_retimer_reg[2][12]  ( .D(\stage_3_output[2][12] ), .CP(clk), 
        .Q(\stage_3_retimer[2][12] ) );
  DFQD1 \stage_3_retimer_reg[2][11]  ( .D(\stage_3_output[2][11] ), .CP(clk), 
        .Q(\stage_3_retimer[2][11] ) );
  DFQD1 \stage_3_retimer_reg[2][10]  ( .D(\stage_3_output[2][10] ), .CP(clk), 
        .Q(\stage_3_retimer[2][10] ) );
  DFQD1 \stage_3_retimer_reg[2][9]  ( .D(\stage_3_output[2][9] ), .CP(clk), 
        .Q(\stage_3_retimer[2][9] ) );
  DFQD1 \stage_3_retimer_reg[2][8]  ( .D(\stage_3_output[2][8] ), .CP(clk), 
        .Q(\stage_3_retimer[2][8] ) );
  DFQD1 \stage_3_retimer_reg[2][7]  ( .D(\stage_3_output[2][7] ), .CP(clk), 
        .Q(\stage_3_retimer[2][7] ) );
  DFQD1 \stage_3_retimer_reg[2][6]  ( .D(\stage_3_output[2][6] ), .CP(clk), 
        .Q(\stage_3_retimer[2][6] ) );
  DFQD1 \stage_3_retimer_reg[2][5]  ( .D(\stage_3_output[2][5] ), .CP(clk), 
        .Q(\stage_3_retimer[2][5] ) );
  DFQD1 \stage_3_retimer_reg[2][4]  ( .D(\stage_3_output[2][4] ), .CP(clk), 
        .Q(\stage_3_retimer[2][4] ) );
  DFQD1 \stage_3_retimer_reg[2][3]  ( .D(\stage_3_output[2][3] ), .CP(clk), 
        .Q(\stage_3_retimer[2][3] ) );
  DFQD1 \stage_3_retimer_reg[2][2]  ( .D(\stage_3_output[2][2] ), .CP(clk), 
        .Q(\stage_3_retimer[2][2] ) );
  DFQD1 \stage_3_retimer_reg[2][1]  ( .D(\stage_3_output[2][1] ), .CP(clk), 
        .Q(\stage_3_retimer[2][1] ) );
  DFQD1 \stage_3_retimer_reg[2][0]  ( .D(\stage_3_output[2][0] ), .CP(clk), 
        .Q(\stage_3_retimer[2][0] ) );
  DFQD1 \stage_3_retimer_reg[1][19]  ( .D(\stage_3_output[1][19] ), .CP(clk), 
        .Q(\stage_3_retimer[1][19] ) );
  DFQD1 \stage_3_retimer_reg[1][18]  ( .D(\stage_3_output[1][18] ), .CP(clk), 
        .Q(\stage_3_retimer[1][18] ) );
  DFQD1 \stage_3_retimer_reg[1][17]  ( .D(\stage_3_output[1][17] ), .CP(clk), 
        .Q(\stage_3_retimer[1][17] ) );
  DFQD1 \stage_3_retimer_reg[1][16]  ( .D(\stage_3_output[1][16] ), .CP(clk), 
        .Q(\stage_3_retimer[1][16] ) );
  DFQD1 \stage_3_retimer_reg[1][15]  ( .D(\stage_3_output[1][15] ), .CP(clk), 
        .Q(\stage_3_retimer[1][15] ) );
  DFQD1 \stage_3_retimer_reg[1][14]  ( .D(\stage_3_output[1][14] ), .CP(clk), 
        .Q(\stage_3_retimer[1][14] ) );
  DFQD1 \stage_3_retimer_reg[1][13]  ( .D(\stage_3_output[1][13] ), .CP(clk), 
        .Q(\stage_3_retimer[1][13] ) );
  DFQD1 \stage_3_retimer_reg[1][12]  ( .D(\stage_3_output[1][12] ), .CP(clk), 
        .Q(\stage_3_retimer[1][12] ) );
  DFQD1 \stage_3_retimer_reg[1][11]  ( .D(\stage_3_output[1][11] ), .CP(clk), 
        .Q(\stage_3_retimer[1][11] ) );
  DFQD1 \stage_3_retimer_reg[1][10]  ( .D(\stage_3_output[1][10] ), .CP(clk), 
        .Q(\stage_3_retimer[1][10] ) );
  DFQD1 \stage_3_retimer_reg[1][9]  ( .D(\stage_3_output[1][9] ), .CP(clk), 
        .Q(\stage_3_retimer[1][9] ) );
  DFQD1 \stage_3_retimer_reg[1][8]  ( .D(\stage_3_output[1][8] ), .CP(clk), 
        .Q(\stage_3_retimer[1][8] ) );
  DFQD1 \stage_3_retimer_reg[1][7]  ( .D(\stage_3_output[1][7] ), .CP(clk), 
        .Q(\stage_3_retimer[1][7] ) );
  DFQD1 \stage_3_retimer_reg[1][6]  ( .D(\stage_3_output[1][6] ), .CP(clk), 
        .Q(\stage_3_retimer[1][6] ) );
  DFQD1 \stage_3_retimer_reg[1][5]  ( .D(\stage_3_output[1][5] ), .CP(clk), 
        .Q(\stage_3_retimer[1][5] ) );
  DFQD1 \stage_3_retimer_reg[1][4]  ( .D(\stage_3_output[1][4] ), .CP(clk), 
        .Q(\stage_3_retimer[1][4] ) );
  DFQD1 \stage_3_retimer_reg[1][3]  ( .D(\stage_3_output[1][3] ), .CP(clk), 
        .Q(\stage_3_retimer[1][3] ) );
  DFQD1 \stage_3_retimer_reg[1][2]  ( .D(\stage_3_output[1][2] ), .CP(clk), 
        .Q(\stage_3_retimer[1][2] ) );
  DFQD1 \stage_3_retimer_reg[1][1]  ( .D(\stage_3_output[1][1] ), .CP(clk), 
        .Q(\stage_3_retimer[1][1] ) );
  DFQD1 \stage_3_retimer_reg[1][0]  ( .D(\stage_3_output[1][0] ), .CP(clk), 
        .Q(\stage_3_retimer[1][0] ) );
  DFQD1 \stage_3_retimer_reg[0][19]  ( .D(\stage_3_output[0][19] ), .CP(clk), 
        .Q(\stage_3_retimer[0][19] ) );
  DFQD1 \stage_3_retimer_reg[0][18]  ( .D(\stage_3_output[0][18] ), .CP(clk), 
        .Q(\stage_3_retimer[0][18] ) );
  DFQD1 \stage_3_retimer_reg[0][17]  ( .D(\stage_3_output[0][17] ), .CP(clk), 
        .Q(\stage_3_retimer[0][17] ) );
  DFQD1 \stage_3_retimer_reg[0][16]  ( .D(\stage_3_output[0][16] ), .CP(clk), 
        .Q(\stage_3_retimer[0][16] ) );
  DFQD1 \stage_3_retimer_reg[0][15]  ( .D(\stage_3_output[0][15] ), .CP(clk), 
        .Q(\stage_3_retimer[0][15] ) );
  DFQD1 \stage_3_retimer_reg[0][14]  ( .D(\stage_3_output[0][14] ), .CP(clk), 
        .Q(\stage_3_retimer[0][14] ) );
  DFQD1 \stage_3_retimer_reg[0][13]  ( .D(\stage_3_output[0][13] ), .CP(clk), 
        .Q(\stage_3_retimer[0][13] ) );
  DFQD1 \stage_3_retimer_reg[0][12]  ( .D(\stage_3_output[0][12] ), .CP(clk), 
        .Q(\stage_3_retimer[0][12] ) );
  DFQD1 \stage_3_retimer_reg[0][11]  ( .D(\stage_3_output[0][11] ), .CP(clk), 
        .Q(\stage_3_retimer[0][11] ) );
  DFQD1 \stage_3_retimer_reg[0][10]  ( .D(\stage_3_output[0][10] ), .CP(clk), 
        .Q(\stage_3_retimer[0][10] ) );
  DFQD1 \stage_3_retimer_reg[0][9]  ( .D(\stage_3_output[0][9] ), .CP(clk), 
        .Q(\stage_3_retimer[0][9] ) );
  DFQD1 \stage_3_retimer_reg[0][8]  ( .D(\stage_3_output[0][8] ), .CP(clk), 
        .Q(\stage_3_retimer[0][8] ) );
  DFQD1 \stage_3_retimer_reg[0][7]  ( .D(\stage_3_output[0][7] ), .CP(clk), 
        .Q(\stage_3_retimer[0][7] ) );
  DFQD1 \stage_3_retimer_reg[0][6]  ( .D(\stage_3_output[0][6] ), .CP(clk), 
        .Q(\stage_3_retimer[0][6] ) );
  DFQD1 \stage_3_retimer_reg[0][5]  ( .D(\stage_3_output[0][5] ), .CP(clk), 
        .Q(\stage_3_retimer[0][5] ) );
  DFQD1 \stage_3_retimer_reg[0][4]  ( .D(\stage_3_output[0][4] ), .CP(clk), 
        .Q(\stage_3_retimer[0][4] ) );
  DFQD1 \stage_3_retimer_reg[0][3]  ( .D(\stage_3_output[0][3] ), .CP(clk), 
        .Q(\stage_3_retimer[0][3] ) );
  DFQD1 \stage_3_retimer_reg[0][2]  ( .D(\stage_3_output[0][2] ), .CP(clk), 
        .Q(\stage_3_retimer[0][2] ) );
  DFQD1 \stage_3_retimer_reg[0][1]  ( .D(\stage_3_output[0][1] ), .CP(clk), 
        .Q(\stage_3_retimer[0][1] ) );
  DFQD1 \stage_3_retimer_reg[0][0]  ( .D(\stage_3_output[0][0] ), .CP(clk), 
        .Q(\stage_3_retimer[0][0] ) );
  DFQD1 \stage_4_retimer_reg[7][19]  ( .D(\stage_4_output[7][19] ), .CP(clk), 
        .Q(out_output[19]) );
  DFQD1 \stage_4_retimer_reg[7][18]  ( .D(\stage_4_output[7][18] ), .CP(clk), 
        .Q(out_output[18]) );
  DFQD1 \stage_4_retimer_reg[7][17]  ( .D(\stage_4_output[7][17] ), .CP(clk), 
        .Q(out_output[17]) );
  DFQD1 \stage_4_retimer_reg[7][16]  ( .D(\stage_4_output[7][16] ), .CP(clk), 
        .Q(out_output[16]) );
  DFQD1 \stage_4_retimer_reg[7][15]  ( .D(\stage_4_output[7][15] ), .CP(clk), 
        .Q(out_output[15]) );
  DFQD1 \stage_4_retimer_reg[7][14]  ( .D(\stage_4_output[7][14] ), .CP(clk), 
        .Q(out_output[14]) );
  DFQD1 \stage_4_retimer_reg[7][13]  ( .D(\stage_4_output[7][13] ), .CP(clk), 
        .Q(out_output[13]) );
  DFQD1 \stage_4_retimer_reg[7][12]  ( .D(\stage_4_output[7][12] ), .CP(clk), 
        .Q(out_output[12]) );
  DFQD1 \stage_4_retimer_reg[7][11]  ( .D(\stage_4_output[7][11] ), .CP(clk), 
        .Q(out_output[11]) );
  DFQD1 \stage_4_retimer_reg[7][10]  ( .D(\stage_4_output[7][10] ), .CP(clk), 
        .Q(out_output[10]) );
  DFQD1 \stage_4_retimer_reg[7][9]  ( .D(\stage_4_output[7][9] ), .CP(clk), 
        .Q(out_output[9]) );
  DFQD1 \stage_4_retimer_reg[7][8]  ( .D(\stage_4_output[7][8] ), .CP(clk), 
        .Q(out_output[8]) );
  DFQD1 \stage_4_retimer_reg[7][7]  ( .D(\stage_4_output[7][7] ), .CP(clk), 
        .Q(out_output[7]) );
  DFQD1 \stage_4_retimer_reg[7][6]  ( .D(\stage_4_output[7][6] ), .CP(clk), 
        .Q(out_output[6]) );
  DFQD1 \stage_4_retimer_reg[7][5]  ( .D(\stage_4_output[7][5] ), .CP(clk), 
        .Q(out_output[5]) );
  DFQD1 \stage_4_retimer_reg[7][4]  ( .D(\stage_4_output[7][4] ), .CP(clk), 
        .Q(out_output[4]) );
  DFQD1 \stage_4_retimer_reg[7][3]  ( .D(\stage_4_output[7][3] ), .CP(clk), 
        .Q(out_output[3]) );
  DFQD1 \stage_4_retimer_reg[7][2]  ( .D(\stage_4_output[7][2] ), .CP(clk), 
        .Q(out_output[2]) );
  DFQD1 \stage_4_retimer_reg[7][1]  ( .D(\stage_4_output[7][1] ), .CP(clk), 
        .Q(out_output[1]) );
  DFQD1 \stage_4_retimer_reg[7][0]  ( .D(\stage_4_output[7][0] ), .CP(clk), 
        .Q(out_output[0]) );
  DFQD1 \stage_4_retimer_reg[6][19]  ( .D(\stage_4_output[6][19] ), .CP(clk), 
        .Q(out_output[39]) );
  DFQD1 \stage_4_retimer_reg[6][18]  ( .D(\stage_4_output[6][18] ), .CP(clk), 
        .Q(out_output[38]) );
  DFQD1 \stage_4_retimer_reg[6][17]  ( .D(\stage_4_output[6][17] ), .CP(clk), 
        .Q(out_output[37]) );
  DFQD1 \stage_4_retimer_reg[6][16]  ( .D(\stage_4_output[6][16] ), .CP(clk), 
        .Q(out_output[36]) );
  DFQD1 \stage_4_retimer_reg[6][15]  ( .D(\stage_4_output[6][15] ), .CP(clk), 
        .Q(out_output[35]) );
  DFQD1 \stage_4_retimer_reg[6][14]  ( .D(\stage_4_output[6][14] ), .CP(clk), 
        .Q(out_output[34]) );
  DFQD1 \stage_4_retimer_reg[6][13]  ( .D(\stage_4_output[6][13] ), .CP(clk), 
        .Q(out_output[33]) );
  DFQD1 \stage_4_retimer_reg[6][12]  ( .D(\stage_4_output[6][12] ), .CP(clk), 
        .Q(out_output[32]) );
  DFQD1 \stage_4_retimer_reg[6][11]  ( .D(\stage_4_output[6][11] ), .CP(clk), 
        .Q(out_output[31]) );
  DFQD1 \stage_4_retimer_reg[6][10]  ( .D(\stage_4_output[6][10] ), .CP(clk), 
        .Q(out_output[30]) );
  DFQD1 \stage_4_retimer_reg[6][9]  ( .D(\stage_4_output[6][9] ), .CP(clk), 
        .Q(out_output[29]) );
  DFQD1 \stage_4_retimer_reg[6][8]  ( .D(\stage_4_output[6][8] ), .CP(clk), 
        .Q(out_output[28]) );
  DFQD1 \stage_4_retimer_reg[6][7]  ( .D(\stage_4_output[6][7] ), .CP(clk), 
        .Q(out_output[27]) );
  DFQD1 \stage_4_retimer_reg[6][6]  ( .D(\stage_4_output[6][6] ), .CP(clk), 
        .Q(out_output[26]) );
  DFQD1 \stage_4_retimer_reg[6][5]  ( .D(\stage_4_output[6][5] ), .CP(clk), 
        .Q(out_output[25]) );
  DFQD1 \stage_4_retimer_reg[6][4]  ( .D(\stage_4_output[6][4] ), .CP(clk), 
        .Q(out_output[24]) );
  DFQD1 \stage_4_retimer_reg[6][3]  ( .D(\stage_4_output[6][3] ), .CP(clk), 
        .Q(out_output[23]) );
  DFQD1 \stage_4_retimer_reg[6][2]  ( .D(\stage_4_output[6][2] ), .CP(clk), 
        .Q(out_output[22]) );
  DFQD1 \stage_4_retimer_reg[6][1]  ( .D(\stage_4_output[6][1] ), .CP(clk), 
        .Q(out_output[21]) );
  DFQD1 \stage_4_retimer_reg[6][0]  ( .D(\stage_4_output[6][0] ), .CP(clk), 
        .Q(out_output[20]) );
  DFQD1 \stage_4_retimer_reg[5][19]  ( .D(\stage_4_output[5][19] ), .CP(clk), 
        .Q(out_output[59]) );
  DFQD1 \stage_4_retimer_reg[5][18]  ( .D(\stage_4_output[5][18] ), .CP(clk), 
        .Q(out_output[58]) );
  DFQD1 \stage_4_retimer_reg[5][17]  ( .D(\stage_4_output[5][17] ), .CP(clk), 
        .Q(out_output[57]) );
  DFQD1 \stage_4_retimer_reg[5][16]  ( .D(\stage_4_output[5][16] ), .CP(clk), 
        .Q(out_output[56]) );
  DFQD1 \stage_4_retimer_reg[5][15]  ( .D(\stage_4_output[5][15] ), .CP(clk), 
        .Q(out_output[55]) );
  DFQD1 \stage_4_retimer_reg[5][14]  ( .D(\stage_4_output[5][14] ), .CP(clk), 
        .Q(out_output[54]) );
  DFQD1 \stage_4_retimer_reg[5][13]  ( .D(\stage_4_output[5][13] ), .CP(clk), 
        .Q(out_output[53]) );
  DFQD1 \stage_4_retimer_reg[5][12]  ( .D(\stage_4_output[5][12] ), .CP(clk), 
        .Q(out_output[52]) );
  DFQD1 \stage_4_retimer_reg[5][11]  ( .D(\stage_4_output[5][11] ), .CP(clk), 
        .Q(out_output[51]) );
  DFQD1 \stage_4_retimer_reg[5][10]  ( .D(\stage_4_output[5][10] ), .CP(clk), 
        .Q(out_output[50]) );
  DFQD1 \stage_4_retimer_reg[5][9]  ( .D(\stage_4_output[5][9] ), .CP(clk), 
        .Q(out_output[49]) );
  DFQD1 \stage_4_retimer_reg[5][8]  ( .D(\stage_4_output[5][8] ), .CP(clk), 
        .Q(out_output[48]) );
  DFQD1 \stage_4_retimer_reg[5][7]  ( .D(\stage_4_output[5][7] ), .CP(clk), 
        .Q(out_output[47]) );
  DFQD1 \stage_4_retimer_reg[5][6]  ( .D(\stage_4_output[5][6] ), .CP(clk), 
        .Q(out_output[46]) );
  DFQD1 \stage_4_retimer_reg[5][5]  ( .D(\stage_4_output[5][5] ), .CP(clk), 
        .Q(out_output[45]) );
  DFQD1 \stage_4_retimer_reg[5][4]  ( .D(\stage_4_output[5][4] ), .CP(clk), 
        .Q(out_output[44]) );
  DFQD1 \stage_4_retimer_reg[5][3]  ( .D(\stage_4_output[5][3] ), .CP(clk), 
        .Q(out_output[43]) );
  DFQD1 \stage_4_retimer_reg[5][2]  ( .D(\stage_4_output[5][2] ), .CP(clk), 
        .Q(out_output[42]) );
  DFQD1 \stage_4_retimer_reg[5][1]  ( .D(\stage_4_output[5][1] ), .CP(clk), 
        .Q(out_output[41]) );
  DFQD1 \stage_4_retimer_reg[5][0]  ( .D(\stage_4_output[5][0] ), .CP(clk), 
        .Q(out_output[40]) );
  DFQD1 \stage_4_retimer_reg[4][19]  ( .D(\stage_4_output[4][19] ), .CP(clk), 
        .Q(out_output[79]) );
  DFQD1 \stage_4_retimer_reg[4][18]  ( .D(\stage_4_output[4][18] ), .CP(clk), 
        .Q(out_output[78]) );
  DFQD1 \stage_4_retimer_reg[4][17]  ( .D(\stage_4_output[4][17] ), .CP(clk), 
        .Q(out_output[77]) );
  DFQD1 \stage_4_retimer_reg[4][16]  ( .D(\stage_4_output[4][16] ), .CP(clk), 
        .Q(out_output[76]) );
  DFQD1 \stage_4_retimer_reg[4][15]  ( .D(\stage_4_output[4][15] ), .CP(clk), 
        .Q(out_output[75]) );
  DFQD1 \stage_4_retimer_reg[4][14]  ( .D(\stage_4_output[4][14] ), .CP(clk), 
        .Q(out_output[74]) );
  DFQD1 \stage_4_retimer_reg[4][13]  ( .D(\stage_4_output[4][13] ), .CP(clk), 
        .Q(out_output[73]) );
  DFQD1 \stage_4_retimer_reg[4][12]  ( .D(\stage_4_output[4][12] ), .CP(clk), 
        .Q(out_output[72]) );
  DFQD1 \stage_4_retimer_reg[4][11]  ( .D(\stage_4_output[4][11] ), .CP(clk), 
        .Q(out_output[71]) );
  DFQD1 \stage_4_retimer_reg[4][10]  ( .D(\stage_4_output[4][10] ), .CP(clk), 
        .Q(out_output[70]) );
  DFQD1 \stage_4_retimer_reg[4][9]  ( .D(\stage_4_output[4][9] ), .CP(clk), 
        .Q(out_output[69]) );
  DFQD1 \stage_4_retimer_reg[4][8]  ( .D(\stage_4_output[4][8] ), .CP(clk), 
        .Q(out_output[68]) );
  DFQD1 \stage_4_retimer_reg[4][7]  ( .D(\stage_4_output[4][7] ), .CP(clk), 
        .Q(out_output[67]) );
  DFQD1 \stage_4_retimer_reg[4][6]  ( .D(\stage_4_output[4][6] ), .CP(clk), 
        .Q(out_output[66]) );
  DFQD1 \stage_4_retimer_reg[4][5]  ( .D(\stage_4_output[4][5] ), .CP(clk), 
        .Q(out_output[65]) );
  DFQD1 \stage_4_retimer_reg[4][4]  ( .D(\stage_4_output[4][4] ), .CP(clk), 
        .Q(out_output[64]) );
  DFQD1 \stage_4_retimer_reg[4][3]  ( .D(\stage_4_output[4][3] ), .CP(clk), 
        .Q(out_output[63]) );
  DFQD1 \stage_4_retimer_reg[4][2]  ( .D(\stage_4_output[4][2] ), .CP(clk), 
        .Q(out_output[62]) );
  DFQD1 \stage_4_retimer_reg[4][1]  ( .D(\stage_4_output[4][1] ), .CP(clk), 
        .Q(out_output[61]) );
  DFQD1 \stage_4_retimer_reg[4][0]  ( .D(\stage_4_output[4][0] ), .CP(clk), 
        .Q(out_output[60]) );
  DFQD1 \stage_4_retimer_reg[3][19]  ( .D(\stage_4_output[3][19] ), .CP(clk), 
        .Q(out_output[99]) );
  DFQD1 \stage_4_retimer_reg[3][18]  ( .D(\stage_4_output[3][18] ), .CP(clk), 
        .Q(out_output[98]) );
  DFQD1 \stage_4_retimer_reg[3][17]  ( .D(\stage_4_output[3][17] ), .CP(clk), 
        .Q(out_output[97]) );
  DFQD1 \stage_4_retimer_reg[3][16]  ( .D(\stage_4_output[3][16] ), .CP(clk), 
        .Q(out_output[96]) );
  DFQD1 \stage_4_retimer_reg[3][15]  ( .D(\stage_4_output[3][15] ), .CP(clk), 
        .Q(out_output[95]) );
  DFQD1 \stage_4_retimer_reg[3][14]  ( .D(\stage_4_output[3][14] ), .CP(clk), 
        .Q(out_output[94]) );
  DFQD1 \stage_4_retimer_reg[3][13]  ( .D(\stage_4_output[3][13] ), .CP(clk), 
        .Q(out_output[93]) );
  DFQD1 \stage_4_retimer_reg[3][12]  ( .D(\stage_4_output[3][12] ), .CP(clk), 
        .Q(out_output[92]) );
  DFQD1 \stage_4_retimer_reg[3][11]  ( .D(\stage_4_output[3][11] ), .CP(clk), 
        .Q(out_output[91]) );
  DFQD1 \stage_4_retimer_reg[3][10]  ( .D(\stage_4_output[3][10] ), .CP(clk), 
        .Q(out_output[90]) );
  DFQD1 \stage_4_retimer_reg[3][9]  ( .D(\stage_4_output[3][9] ), .CP(clk), 
        .Q(out_output[89]) );
  DFQD1 \stage_4_retimer_reg[3][8]  ( .D(\stage_4_output[3][8] ), .CP(clk), 
        .Q(out_output[88]) );
  DFQD1 \stage_4_retimer_reg[3][7]  ( .D(\stage_4_output[3][7] ), .CP(clk), 
        .Q(out_output[87]) );
  DFQD1 \stage_4_retimer_reg[3][6]  ( .D(\stage_4_output[3][6] ), .CP(clk), 
        .Q(out_output[86]) );
  DFQD1 \stage_4_retimer_reg[3][5]  ( .D(\stage_4_output[3][5] ), .CP(clk), 
        .Q(out_output[85]) );
  DFQD1 \stage_4_retimer_reg[3][4]  ( .D(\stage_4_output[3][4] ), .CP(clk), 
        .Q(out_output[84]) );
  DFQD1 \stage_4_retimer_reg[3][3]  ( .D(\stage_4_output[3][3] ), .CP(clk), 
        .Q(out_output[83]) );
  DFQD1 \stage_4_retimer_reg[3][2]  ( .D(\stage_4_output[3][2] ), .CP(clk), 
        .Q(out_output[82]) );
  DFQD1 \stage_4_retimer_reg[3][1]  ( .D(\stage_4_output[3][1] ), .CP(clk), 
        .Q(out_output[81]) );
  DFQD1 \stage_4_retimer_reg[3][0]  ( .D(\stage_4_output[3][0] ), .CP(clk), 
        .Q(out_output[80]) );
  DFQD1 \stage_4_retimer_reg[2][19]  ( .D(\stage_4_output[2][19] ), .CP(clk), 
        .Q(out_output[119]) );
  DFQD1 \stage_4_retimer_reg[2][18]  ( .D(\stage_4_output[2][18] ), .CP(clk), 
        .Q(out_output[118]) );
  DFQD1 \stage_4_retimer_reg[2][17]  ( .D(\stage_4_output[2][17] ), .CP(clk), 
        .Q(out_output[117]) );
  DFQD1 \stage_4_retimer_reg[2][16]  ( .D(\stage_4_output[2][16] ), .CP(clk), 
        .Q(out_output[116]) );
  DFQD1 \stage_4_retimer_reg[2][15]  ( .D(\stage_4_output[2][15] ), .CP(clk), 
        .Q(out_output[115]) );
  DFQD1 \stage_4_retimer_reg[2][14]  ( .D(\stage_4_output[2][14] ), .CP(clk), 
        .Q(out_output[114]) );
  DFQD1 \stage_4_retimer_reg[2][13]  ( .D(\stage_4_output[2][13] ), .CP(clk), 
        .Q(out_output[113]) );
  DFQD1 \stage_4_retimer_reg[2][12]  ( .D(\stage_4_output[2][12] ), .CP(clk), 
        .Q(out_output[112]) );
  DFQD1 \stage_4_retimer_reg[2][11]  ( .D(\stage_4_output[2][11] ), .CP(clk), 
        .Q(out_output[111]) );
  DFQD1 \stage_4_retimer_reg[2][10]  ( .D(\stage_4_output[2][10] ), .CP(clk), 
        .Q(out_output[110]) );
  DFQD1 \stage_4_retimer_reg[2][9]  ( .D(\stage_4_output[2][9] ), .CP(clk), 
        .Q(out_output[109]) );
  DFQD1 \stage_4_retimer_reg[2][8]  ( .D(\stage_4_output[2][8] ), .CP(clk), 
        .Q(out_output[108]) );
  DFQD1 \stage_4_retimer_reg[2][7]  ( .D(\stage_4_output[2][7] ), .CP(clk), 
        .Q(out_output[107]) );
  DFQD1 \stage_4_retimer_reg[2][6]  ( .D(\stage_4_output[2][6] ), .CP(clk), 
        .Q(out_output[106]) );
  DFQD1 \stage_4_retimer_reg[2][5]  ( .D(\stage_4_output[2][5] ), .CP(clk), 
        .Q(out_output[105]) );
  DFQD1 \stage_4_retimer_reg[2][4]  ( .D(\stage_4_output[2][4] ), .CP(clk), 
        .Q(out_output[104]) );
  DFQD1 \stage_4_retimer_reg[2][3]  ( .D(\stage_4_output[2][3] ), .CP(clk), 
        .Q(out_output[103]) );
  DFQD1 \stage_4_retimer_reg[2][2]  ( .D(\stage_4_output[2][2] ), .CP(clk), 
        .Q(out_output[102]) );
  DFQD1 \stage_4_retimer_reg[2][1]  ( .D(\stage_4_output[2][1] ), .CP(clk), 
        .Q(out_output[101]) );
  DFQD1 \stage_4_retimer_reg[2][0]  ( .D(\stage_4_output[2][0] ), .CP(clk), 
        .Q(out_output[100]) );
  DFQD1 \stage_4_retimer_reg[1][19]  ( .D(\stage_4_output[1][19] ), .CP(clk), 
        .Q(out_output[139]) );
  DFQD1 \stage_4_retimer_reg[1][18]  ( .D(\stage_4_output[1][18] ), .CP(clk), 
        .Q(out_output[138]) );
  DFQD1 \stage_4_retimer_reg[1][17]  ( .D(\stage_4_output[1][17] ), .CP(clk), 
        .Q(out_output[137]) );
  DFQD1 \stage_4_retimer_reg[1][16]  ( .D(\stage_4_output[1][16] ), .CP(clk), 
        .Q(out_output[136]) );
  DFQD1 \stage_4_retimer_reg[1][15]  ( .D(\stage_4_output[1][15] ), .CP(clk), 
        .Q(out_output[135]) );
  DFQD1 \stage_4_retimer_reg[1][14]  ( .D(\stage_4_output[1][14] ), .CP(clk), 
        .Q(out_output[134]) );
  DFQD1 \stage_4_retimer_reg[1][13]  ( .D(\stage_4_output[1][13] ), .CP(clk), 
        .Q(out_output[133]) );
  DFQD1 \stage_4_retimer_reg[1][12]  ( .D(\stage_4_output[1][12] ), .CP(clk), 
        .Q(out_output[132]) );
  DFQD1 \stage_4_retimer_reg[1][11]  ( .D(\stage_4_output[1][11] ), .CP(clk), 
        .Q(out_output[131]) );
  DFQD1 \stage_4_retimer_reg[1][10]  ( .D(\stage_4_output[1][10] ), .CP(clk), 
        .Q(out_output[130]) );
  DFQD1 \stage_4_retimer_reg[1][9]  ( .D(\stage_4_output[1][9] ), .CP(clk), 
        .Q(out_output[129]) );
  DFQD1 \stage_4_retimer_reg[1][8]  ( .D(\stage_4_output[1][8] ), .CP(clk), 
        .Q(out_output[128]) );
  DFQD1 \stage_4_retimer_reg[1][7]  ( .D(\stage_4_output[1][7] ), .CP(clk), 
        .Q(out_output[127]) );
  DFQD1 \stage_4_retimer_reg[1][6]  ( .D(\stage_4_output[1][6] ), .CP(clk), 
        .Q(out_output[126]) );
  DFQD1 \stage_4_retimer_reg[1][5]  ( .D(\stage_4_output[1][5] ), .CP(clk), 
        .Q(out_output[125]) );
  DFQD1 \stage_4_retimer_reg[1][4]  ( .D(\stage_4_output[1][4] ), .CP(clk), 
        .Q(out_output[124]) );
  DFQD1 \stage_4_retimer_reg[1][3]  ( .D(\stage_4_output[1][3] ), .CP(clk), 
        .Q(out_output[123]) );
  DFQD1 \stage_4_retimer_reg[1][2]  ( .D(\stage_4_output[1][2] ), .CP(clk), 
        .Q(out_output[122]) );
  DFQD1 \stage_4_retimer_reg[1][1]  ( .D(\stage_4_output[1][1] ), .CP(clk), 
        .Q(out_output[121]) );
  DFQD1 \stage_4_retimer_reg[1][0]  ( .D(\stage_4_output[1][0] ), .CP(clk), 
        .Q(out_output[120]) );
  DFQD1 \stage_4_retimer_reg[0][19]  ( .D(\stage_4_output[0][19] ), .CP(clk), 
        .Q(out_output[159]) );
  DFQD1 \stage_4_retimer_reg[0][18]  ( .D(\stage_4_output[0][18] ), .CP(clk), 
        .Q(out_output[158]) );
  DFQD1 \stage_4_retimer_reg[0][17]  ( .D(\stage_4_output[0][17] ), .CP(clk), 
        .Q(out_output[157]) );
  DFQD1 \stage_4_retimer_reg[0][16]  ( .D(\stage_4_output[0][16] ), .CP(clk), 
        .Q(out_output[156]) );
  DFQD1 \stage_4_retimer_reg[0][15]  ( .D(\stage_4_output[0][15] ), .CP(clk), 
        .Q(out_output[155]) );
  DFQD1 \stage_4_retimer_reg[0][14]  ( .D(\stage_4_output[0][14] ), .CP(clk), 
        .Q(out_output[154]) );
  DFQD1 \stage_4_retimer_reg[0][13]  ( .D(\stage_4_output[0][13] ), .CP(clk), 
        .Q(out_output[153]) );
  DFQD1 \stage_4_retimer_reg[0][12]  ( .D(\stage_4_output[0][12] ), .CP(clk), 
        .Q(out_output[152]) );
  DFQD1 \stage_4_retimer_reg[0][11]  ( .D(\stage_4_output[0][11] ), .CP(clk), 
        .Q(out_output[151]) );
  DFQD1 \stage_4_retimer_reg[0][10]  ( .D(\stage_4_output[0][10] ), .CP(clk), 
        .Q(out_output[150]) );
  DFQD1 \stage_4_retimer_reg[0][9]  ( .D(\stage_4_output[0][9] ), .CP(clk), 
        .Q(out_output[149]) );
  DFQD1 \stage_4_retimer_reg[0][8]  ( .D(\stage_4_output[0][8] ), .CP(clk), 
        .Q(out_output[148]) );
  DFQD1 \stage_4_retimer_reg[0][7]  ( .D(\stage_4_output[0][7] ), .CP(clk), 
        .Q(out_output[147]) );
  DFQD1 \stage_4_retimer_reg[0][6]  ( .D(\stage_4_output[0][6] ), .CP(clk), 
        .Q(out_output[146]) );
  DFQD1 \stage_4_retimer_reg[0][5]  ( .D(\stage_4_output[0][5] ), .CP(clk), 
        .Q(out_output[145]) );
  DFQD1 \stage_4_retimer_reg[0][4]  ( .D(\stage_4_output[0][4] ), .CP(clk), 
        .Q(out_output[144]) );
  DFQD1 \stage_4_retimer_reg[0][3]  ( .D(\stage_4_output[0][3] ), .CP(clk), 
        .Q(out_output[143]) );
  DFQD1 \stage_4_retimer_reg[0][2]  ( .D(\stage_4_output[0][2] ), .CP(clk), 
        .Q(out_output[142]) );
  DFQD1 \stage_4_retimer_reg[0][1]  ( .D(\stage_4_output[0][1] ), .CP(clk), 
        .Q(out_output[141]) );
  DFQD1 \stage_4_retimer_reg[0][0]  ( .D(\stage_4_output[0][0] ), .CP(clk), 
        .Q(out_output[140]) );
  TIEH U3 ( .Z(\*Logic1* ) );
endmodule


module router ( clk, rst, fwd_routing_engine_port_dest, fwd_benes_out_output, 
        fwd_routing_engine_done );
  input [31:0] fwd_routing_engine_port_dest;
  output [159:0] fwd_benes_out_output;
  input clk, rst;
  output fwd_routing_engine_done;
  wire   n2, \output_value[7][15] ;
  wire   [19:0] fwd_routing_engine_control;

  routing_engine_CLOCKED u_fwd_routing_engine ( .port_dest(
        fwd_routing_engine_port_dest), .clk(clk), .rst(rst), .control(
        fwd_routing_engine_control), .done(n2) );
  benes u_fwd_benes ( .in_input({\output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] , 
        \output_value[7][15] , \output_value[7][15] , \output_value[7][15] }), 
        .in_control({\output_value[7][15] , fwd_routing_engine_control[18:16], 
        \output_value[7][15] , fwd_routing_engine_control[14], 
        \output_value[7][15] , fwd_routing_engine_control[12:0]}), .port_en_n(
        {fwd_routing_engine_port_dest[3], fwd_routing_engine_port_dest[7], 
        fwd_routing_engine_port_dest[11], fwd_routing_engine_port_dest[15], 
        fwd_routing_engine_port_dest[19], fwd_routing_engine_port_dest[23], 
        fwd_routing_engine_port_dest[27], fwd_routing_engine_port_dest[31]}), 
        .out_output(fwd_benes_out_output), .clk(\output_value[7][15] ), .rst(
        \output_value[7][15] ) );
  TIEH U1 ( .Z(fwd_routing_engine_done) );
  TIEL U2 ( .ZN(\output_value[7][15] ) );
endmodule

