
module fma_exp_diff_0 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_0 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n604) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n604), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n603) );
  CKXOR2D1 U422 ( .A1(n630), .A2(n603), .Z(n618) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n602) );
  CKXOR2D1 U424 ( .A1(n629), .A2(n602), .Z(n617) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n601) );
  CKXOR2D1 U426 ( .A1(n628), .A2(n601), .Z(n616) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n600) );
  CKXOR2D1 U428 ( .A1(n627), .A2(n600), .Z(n615) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n599) );
  CKXOR2D1 U430 ( .A1(n626), .A2(n599), .Z(n614) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n598) );
  CKXOR2D1 U432 ( .A1(n625), .A2(n598), .Z(n613) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n597) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n597), .Z(n612) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n596) );
  CKXOR2D1 U436 ( .A1(n624), .A2(n596), .Z(n611) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n595) );
  CKXOR2D1 U438 ( .A1(n623), .A2(n595), .Z(n610) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n594) );
  CKXOR2D1 U440 ( .A1(n622), .A2(n594), .Z(n609) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n593) );
  CKXOR2D1 U442 ( .A1(n621), .A2(n593), .Z(n608) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n592) );
  CKXOR2D1 U444 ( .A1(n620), .A2(n592), .Z(n607) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n591) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n590) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n589) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n588) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n587) );
  CKXOR2D1 U450 ( .A1(n619), .A2(n591), .Z(n586) );
  CKXOR2D1 U451 ( .A1(n590), .A2(n589), .Z(n585) );
  CKXOR2D1 U452 ( .A1(n588), .A2(n587), .Z(n584) );
  CKXOR2D1 U453 ( .A1(n586), .A2(n585), .Z(n583) );
  CKXOR2D1 U454 ( .A1(n584), .A2(n583), .Z(n606) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n622) );
  OA21D0 U5 ( .A1(n625), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n625) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n621) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n628), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n620) );
  OAI21D0 U17 ( .A1(n624), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n624) );
  OA31D0 U21 ( .A1(n26), .A2(n627), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n627) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n629), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n619) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n623), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n623)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n626), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n628), .A3(n38), .B(n27), .Z(n626) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n629), .B(N328), .ZN(n628) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n629) );
  CKND0 U56 ( .I(n630), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n630) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n616), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n617), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n618), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n606), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n607), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n608), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n609), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n610), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n611), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n612), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n613), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n614), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n615), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_0 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_0 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_0 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1148, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n1671) );
  CKXOR2D1 U1205 ( .A1(n531), .A2(n1671), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n1680) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n532), .Z(n1670) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n1673), .Z(n1669) );
  CKXOR2D1 U1209 ( .A1(n1670), .A2(n1669), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n1679), .Z(n1678) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n1668) );
  CKXOR2D1 U1212 ( .A1(n1674), .A2(n530), .Z(n1667) );
  CKXOR2D1 U1213 ( .A1(n1668), .A2(n1667), .Z(n1679) );
  CKXOR2D1 U1214 ( .A1(n1676), .A2(n1677), .Z(n1675) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n1666) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n1672), .Z(n1665) );
  CKXOR2D1 U1217 ( .A1(n1666), .A2(n1665), .Z(n1677) );
  fma_lza_0 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_0 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n1148), .SH(exp_diff), .SH_TC(n1148), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n1148) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n1679), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n1676) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n1680), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n1678), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n1679), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n1677), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n1675), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n531), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n1673), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n1673), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n1673) );
  AO21D0 U904 ( .A1(n314), .A2(n1674), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n1674), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n1674) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n531), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n531) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n532), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n532), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n532) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n1672), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n1672) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_0_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_0_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_0 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n23, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_0_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n23), .SH({n77, n76, n74, n75, N11}), .SH_TC(n23), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_0_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n23), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n23) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_0 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_0 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_0 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_0 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n32), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_0 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n32) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_0 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_0 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_7 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_7 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_7 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_7 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_7 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_7 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_7 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_7_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_7_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_7 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_7_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_7_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_7 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_7 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_7 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_7 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_7 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_7 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_7 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_6 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_6 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_6 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_6 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_6 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_6 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_6 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_6_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_6_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_6 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_6_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_6_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_6 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_6 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_6 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_6 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_6 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_6 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_6 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_5 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_5 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_5 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_5 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_5 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_5 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_5 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_5_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_5_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_5 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_5_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_5_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_5 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_5 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_5 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_5 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_5 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_5 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_5 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_4 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_4 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_4 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_4 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_4 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_4 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_4 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_4_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_4_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_4 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_4_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_4_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_4 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_4 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_4 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_4 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_4 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_4 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_4 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_3 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_3 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_3 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_3 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_3 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_3 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_3 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_3_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_3_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_3 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_3_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_3_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_3 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_3 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_3 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_3 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_3 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_3 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_3 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_2 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_2 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_2 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_2 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_2 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_2 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_2 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_2_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_2_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_2 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_2_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_2_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_2 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_2 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_2 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_2 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_2 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_2 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_2 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module fma_exp_diff_1 ( exp_a, exp_b, exp_c, exp_diff_start, fma_byp, exp_diff, 
        exp_ab, exp_ab_greater, exp_ab_less, exp_diff_done );
  input [4:0] exp_a;
  input [4:0] exp_b;
  input [4:0] exp_c;
  output [4:0] exp_diff;
  output [4:0] exp_ab;
  input exp_diff_start, fma_byp;
  output exp_ab_greater, exp_ab_less, exp_diff_done;
  wire   exp_diff_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  assign exp_diff_done = exp_diff_start;

  OAI22D0 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(exp_diff[4]) );
  XNR3D0 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  OAI22D0 U5 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(n7) );
  XNR3D0 U6 ( .A1(n6), .A2(n12), .A3(n13), .ZN(n2) );
  OAI22D0 U7 ( .A1(n14), .A2(n8), .B1(n15), .B2(n16), .ZN(n13) );
  XNR2D0 U8 ( .A1(n17), .A2(n18), .ZN(n6) );
  IND2D0 U9 ( .A1(n19), .B1(n20), .ZN(n18) );
  NR2D0 U10 ( .A1(n12), .A2(n5), .ZN(n17) );
  OAI22D0 U11 ( .A1(n21), .A2(n1), .B1(n4), .B2(n22), .ZN(exp_diff[3]) );
  XNR2D0 U12 ( .A1(n10), .A2(n11), .ZN(n22) );
  XNR2D0 U13 ( .A1(n8), .A2(n9), .ZN(n11) );
  AOI22D0 U14 ( .A1(n23), .A2(exp_c[2]), .B1(n24), .B2(n25), .ZN(n10) );
  XNR2D0 U15 ( .A1(n15), .A2(n16), .ZN(n21) );
  XNR2D0 U16 ( .A1(n8), .A2(n14), .ZN(n16) );
  CKXOR2D0 U17 ( .A1(n20), .A2(n19), .Z(n8) );
  MUX2ND0 U18 ( .I0(n14), .I1(n9), .S(n26), .ZN(n19) );
  NR3D0 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  MAOI22D0 U20 ( .A1(n30), .A2(n23), .B1(n31), .B2(n32), .ZN(n15) );
  OAI22D0 U21 ( .A1(n33), .A2(n1), .B1(n4), .B2(n34), .ZN(exp_diff[2]) );
  XNR2D0 U22 ( .A1(n24), .A2(n25), .ZN(n34) );
  XNR2D0 U23 ( .A1(n23), .A2(n35), .ZN(n25) );
  CKND0 U24 ( .I(n36), .ZN(n24) );
  MAOI222D0 U25 ( .A(exp_c[1]), .B(n37), .C(n38), .ZN(n36) );
  NR2D0 U26 ( .A1(n39), .A2(n40), .ZN(n38) );
  XNR2D0 U27 ( .A1(n31), .A2(n32), .ZN(n33) );
  XNR2D0 U28 ( .A1(n23), .A2(n30), .ZN(n32) );
  XNR2D0 U29 ( .A1(n41), .A2(n28), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n42), .I1(n35), .S(n26), .ZN(n28) );
  NR2D0 U31 ( .A1(n27), .A2(n29), .ZN(n41) );
  MAOI222D0 U32 ( .A(n43), .B(n37), .C(n44), .ZN(n31) );
  XNR2D0 U33 ( .A1(n40), .A2(n29), .ZN(n37) );
  OAI22D0 U34 ( .A1(n1), .A2(n45), .B1(n46), .B2(n4), .ZN(exp_diff[1]) );
  XNR3D0 U35 ( .A1(n47), .A2(exp_c[1]), .A3(n48), .ZN(n46) );
  CKND2D0 U36 ( .A1(n27), .A2(exp_c[0]), .ZN(n47) );
  XNR3D0 U37 ( .A1(n49), .A2(n44), .A3(n48), .ZN(n45) );
  XNR2D0 U38 ( .A1(n27), .A2(n29), .ZN(n48) );
  MUX2ND0 U39 ( .I0(n49), .I1(n50), .S(n26), .ZN(n29) );
  OAI32D0 U40 ( .A1(n1), .A2(n44), .A3(n51), .B1(n4), .B2(n52), .ZN(
        exp_diff[0]) );
  XNR2D0 U41 ( .A1(n40), .A2(n39), .ZN(n52) );
  CKND0 U42 ( .I(exp_ab_less), .ZN(n4) );
  NR2D0 U43 ( .A1(n27), .A2(n53), .ZN(n51) );
  NR2D0 U44 ( .A1(n40), .A2(n54), .ZN(n44) );
  CKND0 U45 ( .I(n27), .ZN(n40) );
  MUX2ND0 U46 ( .I0(n54), .I1(n39), .S(n26), .ZN(n27) );
  INR2D0 U47 ( .A1(n55), .B1(fma_byp), .ZN(exp_ab_less) );
  OAI22D0 U48 ( .A1(n56), .A2(n5), .B1(n57), .B2(n58), .ZN(n55) );
  AOI22D0 U49 ( .A1(n59), .A2(n60), .B1(n14), .B2(exp_c[3]), .ZN(n57) );
  OAI22D0 U50 ( .A1(n35), .A2(n30), .B1(n61), .B2(n62), .ZN(n60) );
  AOI32D0 U51 ( .A1(n54), .A2(n63), .A3(exp_c[0]), .B1(n49), .B2(exp_c[1]), 
        .ZN(n61) );
  CKND0 U52 ( .I(n1), .ZN(exp_ab_greater) );
  IND2D0 U53 ( .A1(fma_byp), .B1(n26), .ZN(n1) );
  OAI22D0 U54 ( .A1(exp_c[4]), .A2(n12), .B1(n64), .B2(n58), .ZN(n26) );
  XNR2D0 U55 ( .A1(n56), .A2(n5), .ZN(n58) );
  CKND0 U56 ( .I(exp_c[4]), .ZN(n5) );
  AOI22D0 U57 ( .A1(n59), .A2(n65), .B1(n66), .B2(n9), .ZN(n64) );
  OAI22D0 U58 ( .A1(exp_c[2]), .A2(n42), .B1(n67), .B2(n62), .ZN(n65) );
  XNR2D0 U59 ( .A1(n30), .A2(n35), .ZN(n62) );
  CKND0 U60 ( .I(exp_c[2]), .ZN(n35) );
  AOI32D0 U61 ( .A1(n53), .A2(n39), .A3(n63), .B1(n43), .B2(n50), .ZN(n67) );
  XNR2D0 U62 ( .A1(n49), .A2(n50), .ZN(n63) );
  CKND0 U63 ( .I(exp_c[1]), .ZN(n50) );
  CKND0 U64 ( .I(exp_c[0]), .ZN(n39) );
  XNR2D0 U65 ( .A1(n14), .A2(n9), .ZN(n59) );
  CKND0 U66 ( .I(exp_c[3]), .ZN(n9) );
  NR2D0 U67 ( .A1(fma_byp), .A2(n12), .ZN(exp_ab[4]) );
  CKND0 U68 ( .I(n56), .ZN(n12) );
  CKND2D0 U69 ( .A1(n68), .A2(n69), .ZN(n56) );
  NR2D0 U70 ( .A1(fma_byp), .A2(n14), .ZN(exp_ab[3]) );
  CKND0 U71 ( .I(n66), .ZN(n14) );
  CKND2D0 U72 ( .A1(n70), .A2(n71), .ZN(n66) );
  XNR2D0 U73 ( .A1(n72), .A2(n73), .ZN(n71) );
  NR2D0 U74 ( .A1(fma_byp), .A2(n42), .ZN(exp_ab[2]) );
  CKND0 U75 ( .I(n30), .ZN(n42) );
  CKND2D0 U76 ( .A1(n74), .A2(n70), .ZN(n30) );
  XNR2D0 U77 ( .A1(n75), .A2(n76), .ZN(n74) );
  NR2D0 U78 ( .A1(fma_byp), .A2(n49), .ZN(exp_ab[1]) );
  CKND0 U79 ( .I(n43), .ZN(n49) );
  CKND2D0 U80 ( .A1(n77), .A2(n70), .ZN(n43) );
  XNR3D0 U81 ( .A1(exp_b[1]), .A2(exp_a[1]), .A3(n78), .ZN(n77) );
  NR2D0 U82 ( .A1(fma_byp), .A2(n54), .ZN(exp_ab[0]) );
  CKND0 U83 ( .I(n53), .ZN(n54) );
  OAI21D0 U84 ( .A1(n79), .A2(n78), .B(n70), .ZN(n53) );
  MAOI22D0 U85 ( .A1(exp_b[4]), .A2(exp_a[4]), .B1(n68), .B2(n69), .ZN(n70) );
  NR2D0 U86 ( .A1(exp_a[4]), .A2(exp_b[4]), .ZN(n69) );
  OA21D0 U87 ( .A1(n72), .A2(n73), .B(n80), .Z(n68) );
  OAI21D0 U88 ( .A1(exp_b[3]), .A2(exp_a[3]), .B(n80), .ZN(n73) );
  CKND2D0 U89 ( .A1(exp_b[3]), .A2(exp_a[3]), .ZN(n80) );
  OA21D0 U90 ( .A1(n75), .A2(n76), .B(n81), .Z(n72) );
  MAOI222D0 U91 ( .A(exp_b[1]), .B(n78), .C(exp_a[1]), .ZN(n76) );
  OAI21D0 U92 ( .A1(exp_b[2]), .A2(exp_a[2]), .B(n81), .ZN(n75) );
  CKND2D0 U93 ( .A1(exp_b[2]), .A2(exp_a[2]), .ZN(n81) );
  AN2D0 U94 ( .A1(exp_b[0]), .A2(exp_a[0]), .Z(n78) );
  NR2D0 U95 ( .A1(exp_b[0]), .A2(exp_a[0]), .ZN(n79) );
endmodule


module fma_mult_tree_1 ( mantissa_a, mantissa_b, sign_a, sign_b, fma_byp, 
        a_equals_one, b_equals_one, mult_start, mantissa_ab, sign_ab, 
        mult_done );
  input [9:0] mantissa_a;
  input [9:0] mantissa_b;
  output [19:0] mantissa_ab;
  input sign_a, sign_b, fma_byp, a_equals_one, b_equals_one, mult_start;
  output sign_ab, mult_done;
  wire   mult_start, N37, N66, N93, N118, N141, N142, N251, N255, N317, N323,
         N324, N325, N326, N327, N328, N329, N332, N333, N336, N337, N340,
         N341, N344, N345, N348, N349, N352, N353, N356, N357, N360, N361,
         N364, N365, N368, N369, N373, N470, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541;
  assign mult_done = mult_start;

  CKXOR2D1 U419 ( .A1(N373), .A2(N323), .Z(n520) );
  CKXOR2D1 U420 ( .A1(N324), .A2(n520), .Z(N470) );
  CKXOR2D1 U421 ( .A1(N325), .A2(N326), .Z(n521) );
  CKXOR2D1 U422 ( .A1(n495), .A2(n521), .Z(n507) );
  CKXOR2D1 U423 ( .A1(N327), .A2(N328), .Z(n522) );
  CKXOR2D1 U424 ( .A1(n496), .A2(n522), .Z(n508) );
  CKXOR2D1 U425 ( .A1(N329), .A2(N332), .Z(n523) );
  CKXOR2D1 U426 ( .A1(n497), .A2(n523), .Z(n509) );
  CKXOR2D1 U427 ( .A1(N333), .A2(N336), .Z(n524) );
  CKXOR2D1 U428 ( .A1(n498), .A2(n524), .Z(n510) );
  CKXOR2D1 U429 ( .A1(N337), .A2(N340), .Z(n525) );
  CKXOR2D1 U430 ( .A1(n499), .A2(n525), .Z(n511) );
  CKXOR2D1 U431 ( .A1(N341), .A2(N344), .Z(n526) );
  CKXOR2D1 U432 ( .A1(n500), .A2(n526), .Z(n512) );
  CKXOR2D1 U433 ( .A1(N345), .A2(N348), .Z(n527) );
  CKXOR2D1 U434 ( .A1(n494), .A2(n527), .Z(n513) );
  CKXOR2D1 U435 ( .A1(N349), .A2(N352), .Z(n528) );
  CKXOR2D1 U436 ( .A1(n501), .A2(n528), .Z(n514) );
  CKXOR2D1 U437 ( .A1(N353), .A2(N356), .Z(n529) );
  CKXOR2D1 U438 ( .A1(n502), .A2(n529), .Z(n515) );
  CKXOR2D1 U439 ( .A1(N357), .A2(N360), .Z(n530) );
  CKXOR2D1 U440 ( .A1(n503), .A2(n530), .Z(n516) );
  CKXOR2D1 U441 ( .A1(N361), .A2(N364), .Z(n531) );
  CKXOR2D1 U442 ( .A1(n504), .A2(n531), .Z(n517) );
  CKXOR2D1 U443 ( .A1(N365), .A2(N368), .Z(n532) );
  CKXOR2D1 U444 ( .A1(n505), .A2(n532), .Z(n518) );
  CKXOR2D1 U445 ( .A1(N142), .A2(N37), .Z(n533) );
  CKXOR2D1 U446 ( .A1(N66), .A2(N93), .Z(n534) );
  CKXOR2D1 U447 ( .A1(N118), .A2(N141), .Z(n535) );
  CKXOR2D1 U448 ( .A1(N251), .A2(N255), .Z(n536) );
  CKXOR2D1 U449 ( .A1(N317), .A2(N369), .Z(n537) );
  CKXOR2D1 U450 ( .A1(n506), .A2(n533), .Z(n538) );
  CKXOR2D1 U451 ( .A1(n534), .A2(n535), .Z(n539) );
  CKXOR2D1 U452 ( .A1(n536), .A2(n537), .Z(n540) );
  CKXOR2D1 U453 ( .A1(n538), .A2(n539), .Z(n541) );
  CKXOR2D1 U454 ( .A1(n540), .A2(n541), .Z(n519) );
  CKXOR2D0 U2 ( .A1(sign_b), .A2(sign_a), .Z(sign_ab) );
  CKND0 U3 ( .I(n1), .ZN(n494) );
  OA211D0 U4 ( .A1(n2), .A2(n3), .B(n4), .C(n5), .Z(n503) );
  OA21D0 U5 ( .A1(n500), .A2(n6), .B(n7), .Z(n3) );
  OA221D0 U6 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C(n12), .Z(n500) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(n9) );
  AOI21D0 U8 ( .A1(n15), .A2(n16), .B(n17), .ZN(n504) );
  MOAI22D0 U9 ( .A1(n18), .A2(n5), .B1(N357), .B2(N360), .ZN(n17) );
  OAI21D0 U10 ( .A1(n19), .A2(n2), .B(n4), .ZN(n16) );
  AOI21D0 U11 ( .A1(n1), .A2(n20), .B(n21), .ZN(n19) );
  OAI22D0 U12 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(n1) );
  OA221D0 U13 ( .A1(n26), .A2(n27), .B1(n10), .B2(n497), .C(n28), .Z(n24) );
  ND3D0 U14 ( .A1(N332), .A2(n14), .A3(n13), .ZN(n10) );
  CKND0 U15 ( .I(n18), .ZN(n15) );
  AOI21D0 U16 ( .A1(n29), .A2(n30), .B(n31), .ZN(n505) );
  OAI21D0 U17 ( .A1(n501), .A2(n2), .B(n4), .ZN(n30) );
  CKND2D0 U18 ( .A1(n32), .A2(n33), .ZN(n4) );
  OAI21D0 U19 ( .A1(N349), .A2(N352), .B(n33), .ZN(n2) );
  IAO21D0 U20 ( .A1(n34), .A2(n6), .B(n35), .ZN(n501) );
  OA31D0 U21 ( .A1(n26), .A2(n498), .A3(n36), .B(n12), .Z(n34) );
  AOI31D0 U22 ( .A1(N336), .A2(N333), .A3(n14), .B(n37), .ZN(n12) );
  CKND0 U23 ( .I(n28), .ZN(n37) );
  CKND0 U24 ( .I(n26), .ZN(n14) );
  OA21D0 U25 ( .A1(n38), .A2(n11), .B(n8), .Z(n498) );
  CKND2D0 U26 ( .A1(N332), .A2(n39), .ZN(n8) );
  OAI21D0 U27 ( .A1(n40), .A2(n41), .B(n42), .ZN(n39) );
  OR2D0 U28 ( .A1(n496), .A2(n40), .Z(n11) );
  CKND0 U29 ( .I(N328), .ZN(n40) );
  CKND0 U30 ( .I(n43), .ZN(n506) );
  MAOI222D0 U31 ( .A(n44), .B(n45), .C(n46), .ZN(n43) );
  MAOI22D0 U32 ( .A1(n47), .A2(n48), .B1(n49), .B2(n50), .ZN(n46) );
  CKXOR2D0 U33 ( .A1(n51), .A2(n52), .Z(n45) );
  CKND0 U34 ( .I(n53), .ZN(n52) );
  AOI31D0 U35 ( .A1(n33), .A2(n54), .A3(n29), .B(n31), .ZN(n44) );
  MAOI222D0 U36 ( .A(n55), .B(n56), .C(n57), .ZN(n31) );
  AOI22D0 U37 ( .A1(n58), .A2(n59), .B1(n60), .B2(n61), .ZN(n57) );
  MAOI22D0 U38 ( .A1(N360), .A2(N357), .B1(n5), .B2(n18), .ZN(n56) );
  CKND2D0 U39 ( .A1(N356), .A2(N353), .ZN(n5) );
  IAO21D0 U40 ( .A1(N361), .A2(N364), .B(n18), .ZN(n29) );
  XNR2D0 U41 ( .A1(N360), .A2(N357), .ZN(n18) );
  CKND0 U42 ( .I(n502), .ZN(n54) );
  OAI32D0 U43 ( .A1(n62), .A2(n32), .A3(n35), .B1(N349), .B2(N352), .ZN(n502)
         );
  CKND0 U44 ( .I(n7), .ZN(n35) );
  AOI31D0 U45 ( .A1(N344), .A2(n20), .A3(N341), .B(n21), .ZN(n7) );
  AN2D0 U46 ( .A1(N348), .A2(N345), .Z(n21) );
  CKND0 U47 ( .I(n63), .ZN(n20) );
  AN2D0 U48 ( .A1(N352), .A2(N349), .Z(n32) );
  OAI33D0 U49 ( .A1(n28), .A2(n63), .A3(n25), .B1(n6), .B2(n499), .B3(n26), 
        .ZN(n62) );
  NR2D0 U50 ( .A1(N340), .A2(N337), .ZN(n26) );
  OA31D0 U51 ( .A1(n36), .A2(n497), .A3(n38), .B(n27), .Z(n499) );
  AOI32D0 U52 ( .A1(N329), .A2(N332), .A3(n13), .B1(N333), .B2(N336), .ZN(n27)
         );
  CKND0 U53 ( .I(n36), .ZN(n13) );
  IOA21D0 U54 ( .A1(n41), .A2(n496), .B(N328), .ZN(n497) );
  OAI21D0 U55 ( .A1(N325), .A2(n64), .B(N326), .ZN(n496) );
  CKND0 U56 ( .I(n495), .ZN(n64) );
  OAI21D0 U57 ( .A1(N373), .A2(N323), .B(N324), .ZN(n495) );
  XNR2D0 U58 ( .A1(N336), .A2(N333), .ZN(n36) );
  OR2D0 U59 ( .A1(n25), .A2(n63), .Z(n6) );
  CKXOR2D0 U60 ( .A1(N344), .A2(n22), .Z(n25) );
  CKND0 U61 ( .I(N341), .ZN(n22) );
  NR2D0 U62 ( .A1(N348), .A2(N345), .ZN(n63) );
  CKND2D0 U63 ( .A1(N340), .A2(N337), .ZN(n28) );
  CKXOR2D0 U64 ( .A1(N353), .A2(N356), .Z(n33) );
  OAI222D0 U65 ( .A1(n509), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(mantissa_ab[9]) );
  OAI222D0 U66 ( .A1(n508), .A2(n65), .B1(n70), .B2(n67), .C1(n71), .C2(n69), 
        .ZN(mantissa_ab[8]) );
  OAI222D0 U67 ( .A1(n507), .A2(n65), .B1(n72), .B2(n67), .C1(n73), .C2(n69), 
        .ZN(mantissa_ab[7]) );
  CKND0 U68 ( .I(mantissa_a[7]), .ZN(n72) );
  AO222D0 U69 ( .A1(N470), .A2(n74), .B1(n75), .B2(mantissa_a[6]), .C1(n76), 
        .C2(mantissa_b[6]), .Z(mantissa_ab[6]) );
  CKND0 U70 ( .I(n69), .ZN(n76) );
  OAI222D0 U71 ( .A1(n77), .A2(n67), .B1(n78), .B2(n65), .C1(n79), .C2(n69), 
        .ZN(mantissa_ab[5]) );
  CKXOR2D0 U72 ( .A1(n80), .A2(n81), .Z(n78) );
  CKND0 U73 ( .I(mantissa_a[5]), .ZN(n77) );
  OAI222D0 U74 ( .A1(n82), .A2(n67), .B1(n83), .B2(n65), .C1(n84), .C2(n69), 
        .ZN(mantissa_ab[4]) );
  XNR2D0 U75 ( .A1(n85), .A2(n86), .ZN(n83) );
  CKND0 U76 ( .I(mantissa_a[4]), .ZN(n82) );
  OAI222D0 U77 ( .A1(n87), .A2(n67), .B1(n88), .B2(n65), .C1(n89), .C2(n69), 
        .ZN(mantissa_ab[3]) );
  CKXOR2D0 U78 ( .A1(n90), .A2(n91), .Z(n88) );
  CKND0 U79 ( .I(mantissa_a[3]), .ZN(n87) );
  OAI222D0 U80 ( .A1(n92), .A2(n67), .B1(n65), .B2(n93), .C1(n94), .C2(n69), 
        .ZN(mantissa_ab[2]) );
  XNR2D0 U81 ( .A1(n95), .A2(n96), .ZN(n93) );
  CKND0 U82 ( .I(mantissa_a[2]), .ZN(n92) );
  OAI222D0 U83 ( .A1(n97), .A2(n67), .B1(n65), .B2(n98), .C1(n99), .C2(n69), 
        .ZN(mantissa_ab[1]) );
  CKXOR2D0 U84 ( .A1(n100), .A2(n101), .Z(n98) );
  CKND0 U85 ( .I(mantissa_a[1]), .ZN(n97) );
  NR2D0 U86 ( .A1(n519), .A2(n65), .ZN(mantissa_ab[19]) );
  NR2D0 U87 ( .A1(n518), .A2(n65), .ZN(mantissa_ab[18]) );
  NR2D0 U88 ( .A1(n517), .A2(n65), .ZN(mantissa_ab[17]) );
  NR2D0 U89 ( .A1(n516), .A2(n65), .ZN(mantissa_ab[16]) );
  NR2D0 U90 ( .A1(n515), .A2(n65), .ZN(mantissa_ab[15]) );
  NR2D0 U91 ( .A1(n514), .A2(n65), .ZN(mantissa_ab[14]) );
  NR2D0 U92 ( .A1(n513), .A2(n65), .ZN(mantissa_ab[13]) );
  NR2D0 U93 ( .A1(n512), .A2(n65), .ZN(mantissa_ab[12]) );
  NR2D0 U94 ( .A1(n511), .A2(n65), .ZN(mantissa_ab[11]) );
  NR2D0 U95 ( .A1(n510), .A2(n65), .ZN(mantissa_ab[10]) );
  OAI222D0 U96 ( .A1(n102), .A2(n67), .B1(n65), .B2(n103), .C1(n104), .C2(n69), 
        .ZN(mantissa_ab[0]) );
  IND2D0 U97 ( .A1(fma_byp), .B1(a_equals_one), .ZN(n69) );
  CKXOR2D0 U98 ( .A1(n105), .A2(n99), .Z(n103) );
  CKND0 U99 ( .I(n74), .ZN(n65) );
  CKND0 U100 ( .I(n75), .ZN(n67) );
  NR3D0 U101 ( .A1(a_equals_one), .A2(fma_byp), .A3(n74), .ZN(n75) );
  NR3D0 U102 ( .A1(fma_byp), .A2(b_equals_one), .A3(a_equals_one), .ZN(n74) );
  CKND0 U103 ( .I(n106), .ZN(N93) );
  CKND0 U104 ( .I(n107), .ZN(N66) );
  INR2D0 U105 ( .A1(n80), .B1(n81), .ZN(N373) );
  CKND2D0 U106 ( .A1(n86), .A2(n85), .ZN(n81) );
  XNR2D0 U107 ( .A1(n108), .A2(n109), .ZN(n85) );
  CKND2D0 U108 ( .A1(n110), .A2(n111), .ZN(n109) );
  INR2D0 U109 ( .A1(n90), .B1(n91), .ZN(n86) );
  CKND2D0 U110 ( .A1(n95), .A2(n96), .ZN(n91) );
  CKXOR2D0 U111 ( .A1(n112), .A2(n89), .Z(n96) );
  CKXOR2D0 U112 ( .A1(n113), .A2(n114), .Z(n95) );
  CKXOR2D0 U113 ( .A1(n110), .A2(n111), .Z(n90) );
  XNR2D0 U114 ( .A1(n115), .A2(n116), .ZN(n80) );
  MOAI22D0 U115 ( .A1(n117), .A2(n118), .B1(n53), .B2(n51), .ZN(N369) );
  CKXOR2D0 U116 ( .A1(n51), .A2(n53), .Z(N368) );
  CKXOR2D0 U117 ( .A1(n119), .A2(n120), .Z(n53) );
  CKXOR2D0 U118 ( .A1(n117), .A2(n118), .Z(n51) );
  OA21D0 U119 ( .A1(n121), .A2(n122), .B(n123), .Z(n118) );
  AN2D0 U120 ( .A1(n124), .A2(n125), .Z(n117) );
  MOAI22D0 U121 ( .A1(n50), .A2(n49), .B1(n48), .B2(n47), .ZN(N365) );
  CKND0 U122 ( .I(n55), .ZN(N364) );
  XNR2D0 U123 ( .A1(n50), .A2(n49), .ZN(n55) );
  OAI21D0 U124 ( .A1(n142), .A2(n126), .B(n124), .ZN(n49) );
  CKND2D0 U125 ( .A1(n142), .A2(n126), .ZN(n124) );
  OA21D0 U126 ( .A1(n127), .A2(N251), .B(n125), .Z(n126) );
  CKND2D0 U127 ( .A1(n127), .A2(N251), .ZN(n125) );
  OA21D0 U128 ( .A1(n128), .A2(n129), .B(n123), .Z(n127) );
  CKND2D0 U129 ( .A1(n128), .A2(n129), .ZN(n123) );
  IAO21D0 U130 ( .A1(n130), .A2(n131), .B(n73), .ZN(n129) );
  CKXOR2D0 U131 ( .A1(n121), .A2(n122), .Z(n128) );
  CKND2D0 U132 ( .A1(mantissa_b[9]), .A2(mantissa_a[7]), .ZN(n122) );
  CKXOR2D0 U133 ( .A1(n132), .A2(n133), .Z(n121) );
  CKND2D0 U134 ( .A1(n134), .A2(n135), .ZN(n133) );
  XNR2D0 U135 ( .A1(n48), .A2(n47), .ZN(n50) );
  OAI21D0 U136 ( .A1(n136), .A2(n137), .B(n138), .ZN(n47) );
  CKND2D0 U137 ( .A1(n139), .A2(n140), .ZN(n48) );
  AO22D0 U138 ( .A1(n59), .A2(n58), .B1(n61), .B2(n60), .Z(N361) );
  CKXOR2D0 U139 ( .A1(n59), .A2(n58), .Z(N360) );
  OA21D0 U140 ( .A1(n141), .A2(n142), .B(n139), .Z(n58) );
  CKND2D0 U141 ( .A1(n141), .A2(n142), .ZN(n139) );
  OA21D0 U142 ( .A1(n143), .A2(N251), .B(n140), .Z(n141) );
  CKND2D0 U143 ( .A1(n143), .A2(N251), .ZN(n140) );
  OA21D0 U144 ( .A1(n144), .A2(n145), .B(n138), .Z(n143) );
  CKND2D0 U145 ( .A1(n144), .A2(n145), .ZN(n138) );
  CKXOR2D0 U146 ( .A1(n131), .A2(n130), .Z(n145) );
  CKXOR2D0 U147 ( .A1(n136), .A2(n137), .Z(n144) );
  CKND2D0 U148 ( .A1(mantissa_b[9]), .A2(mantissa_a[6]), .ZN(n137) );
  XNR2D0 U149 ( .A1(n134), .A2(n135), .ZN(n136) );
  CKXOR2D0 U150 ( .A1(n61), .A2(n60), .Z(n59) );
  OAI21D0 U151 ( .A1(n146), .A2(n147), .B(n148), .ZN(n60) );
  CKND2D0 U152 ( .A1(n149), .A2(n150), .ZN(n61) );
  OAI22D0 U153 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .ZN(N357) );
  CKXOR2D0 U154 ( .A1(n153), .A2(n154), .Z(N356) );
  OAI21D0 U155 ( .A1(n155), .A2(n142), .B(n149), .ZN(n154) );
  CKND2D0 U156 ( .A1(n155), .A2(n142), .ZN(n149) );
  OA21D0 U157 ( .A1(N37), .A2(n156), .B(n157), .Z(n142) );
  OA21D0 U158 ( .A1(n158), .A2(n159), .B(n150), .Z(n155) );
  CKND2D0 U159 ( .A1(n158), .A2(n159), .ZN(n150) );
  OAI21D0 U160 ( .A1(n107), .A2(n160), .B(n161), .ZN(n159) );
  OA21D0 U161 ( .A1(n162), .A2(n163), .B(n148), .Z(n158) );
  CKND2D0 U162 ( .A1(n162), .A2(n163), .ZN(n148) );
  XNR2D0 U163 ( .A1(n164), .A2(n165), .ZN(n163) );
  CKND2D0 U164 ( .A1(n166), .A2(n167), .ZN(n165) );
  CKXOR2D0 U165 ( .A1(n146), .A2(n147), .Z(n162) );
  CKND2D0 U166 ( .A1(mantissa_b[9]), .A2(mantissa_a[5]), .ZN(n147) );
  XNR2D0 U167 ( .A1(n168), .A2(n169), .ZN(n146) );
  AN2D0 U168 ( .A1(n170), .A2(n171), .Z(n168) );
  XNR2D0 U169 ( .A1(n151), .A2(n152), .ZN(n153) );
  OA21D0 U170 ( .A1(n172), .A2(n173), .B(n174), .Z(n152) );
  AN2D0 U171 ( .A1(n175), .A2(n176), .Z(n151) );
  OAI22D0 U172 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .ZN(N353) );
  CKXOR2D0 U173 ( .A1(n179), .A2(n180), .Z(N352) );
  OAI21D0 U174 ( .A1(n181), .A2(n182), .B(n175), .ZN(n180) );
  CKND2D0 U175 ( .A1(n181), .A2(n182), .ZN(n175) );
  OA21D0 U176 ( .A1(N37), .A2(n183), .B(n161), .Z(n182) );
  CKND2D0 U177 ( .A1(n183), .A2(N37), .ZN(n161) );
  CKXOR2D0 U178 ( .A1(n107), .A2(n160), .Z(n183) );
  XNR2D0 U179 ( .A1(n184), .A2(n185), .ZN(n160) );
  OA21D0 U180 ( .A1(n186), .A2(n187), .B(n176), .Z(n181) );
  CKND2D0 U181 ( .A1(n186), .A2(n187), .ZN(n176) );
  OAI21D0 U182 ( .A1(n107), .A2(n188), .B(n189), .ZN(n187) );
  OA21D0 U183 ( .A1(n190), .A2(n191), .B(n174), .Z(n186) );
  CKND2D0 U184 ( .A1(n190), .A2(n191), .ZN(n174) );
  CKXOR2D0 U185 ( .A1(n166), .A2(n167), .Z(n191) );
  CKXOR2D0 U186 ( .A1(n172), .A2(n173), .Z(n190) );
  CKND2D0 U187 ( .A1(mantissa_b[9]), .A2(mantissa_a[4]), .ZN(n173) );
  CKXOR2D0 U188 ( .A1(n192), .A2(n170), .Z(n172) );
  XNR2D0 U189 ( .A1(n177), .A2(n178), .ZN(n179) );
  OA21D0 U190 ( .A1(n193), .A2(n194), .B(n195), .Z(n178) );
  AN2D0 U191 ( .A1(n196), .A2(n197), .Z(n177) );
  OAI22D0 U192 ( .A1(n198), .A2(n199), .B1(n200), .B2(n201), .ZN(N349) );
  CKXOR2D0 U193 ( .A1(n200), .A2(n201), .Z(N348) );
  OAI21D0 U194 ( .A1(n202), .A2(n203), .B(n196), .ZN(n201) );
  CKND2D0 U195 ( .A1(n202), .A2(n203), .ZN(n196) );
  OA21D0 U196 ( .A1(N37), .A2(n204), .B(n189), .Z(n203) );
  CKND2D0 U197 ( .A1(n204), .A2(N37), .ZN(n189) );
  CKXOR2D0 U198 ( .A1(n107), .A2(n188), .Z(n204) );
  CKXOR2D0 U199 ( .A1(n205), .A2(n206), .Z(n188) );
  CKND2D0 U200 ( .A1(n207), .A2(n208), .ZN(n206) );
  OA21D0 U201 ( .A1(n209), .A2(n210), .B(n197), .Z(n202) );
  CKND2D0 U202 ( .A1(n209), .A2(n210), .ZN(n197) );
  OAI21D0 U203 ( .A1(n211), .A2(n212), .B(n213), .ZN(n210) );
  OA21D0 U204 ( .A1(n214), .A2(n215), .B(n195), .Z(n209) );
  CKND2D0 U205 ( .A1(n214), .A2(n215), .ZN(n195) );
  CKXOR2D0 U206 ( .A1(n216), .A2(n217), .Z(n215) );
  NR2D0 U207 ( .A1(n218), .A2(n219), .ZN(n216) );
  CKXOR2D0 U208 ( .A1(n193), .A2(n194), .Z(n214) );
  CKND2D0 U209 ( .A1(mantissa_b[9]), .A2(mantissa_a[3]), .ZN(n194) );
  XNR2D0 U210 ( .A1(n220), .A2(n221), .ZN(n193) );
  CKND2D0 U211 ( .A1(n222), .A2(n223), .ZN(n221) );
  XNR2D0 U212 ( .A1(n198), .A2(n199), .ZN(n200) );
  OA21D0 U213 ( .A1(n224), .A2(n225), .B(n226), .Z(n199) );
  AN2D0 U214 ( .A1(n227), .A2(n228), .Z(n198) );
  OAI22D0 U215 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(N345) );
  CKND0 U216 ( .I(n23), .ZN(N344) );
  XNR2D0 U217 ( .A1(n231), .A2(n232), .ZN(n23) );
  OAI21D0 U218 ( .A1(n233), .A2(n234), .B(n227), .ZN(n232) );
  CKND2D0 U219 ( .A1(n233), .A2(n234), .ZN(n227) );
  OA21D0 U220 ( .A1(N37), .A2(n235), .B(n213), .Z(n234) );
  CKND2D0 U221 ( .A1(n235), .A2(N37), .ZN(n213) );
  CKXOR2D0 U222 ( .A1(n211), .A2(n212), .Z(n235) );
  XNR2D0 U223 ( .A1(n207), .A2(n208), .ZN(n212) );
  XNR2D0 U224 ( .A1(n236), .A2(n237), .ZN(n211) );
  OA21D0 U225 ( .A1(n238), .A2(n239), .B(n228), .Z(n233) );
  CKND2D0 U226 ( .A1(n238), .A2(n239), .ZN(n228) );
  OAI21D0 U227 ( .A1(n240), .A2(n241), .B(n242), .ZN(n239) );
  OA21D0 U228 ( .A1(n243), .A2(n244), .B(n226), .Z(n238) );
  CKND2D0 U229 ( .A1(n243), .A2(n244), .ZN(n226) );
  CKXOR2D0 U230 ( .A1(n219), .A2(n218), .Z(n244) );
  CKXOR2D0 U231 ( .A1(n224), .A2(n225), .Z(n243) );
  CKND2D0 U232 ( .A1(mantissa_b[9]), .A2(mantissa_a[2]), .ZN(n225) );
  XNR2D0 U233 ( .A1(n222), .A2(n223), .ZN(n224) );
  XNR2D0 U234 ( .A1(n229), .A2(n230), .ZN(n231) );
  OA21D0 U235 ( .A1(n245), .A2(n246), .B(n247), .Z(n230) );
  AN2D0 U236 ( .A1(n248), .A2(n249), .Z(n229) );
  OAI22D0 U237 ( .A1(n250), .A2(n251), .B1(n252), .B2(n253), .ZN(N341) );
  CKXOR2D0 U238 ( .A1(n252), .A2(n253), .Z(N340) );
  OAI21D0 U239 ( .A1(n254), .A2(n255), .B(n248), .ZN(n253) );
  CKND2D0 U240 ( .A1(n254), .A2(n255), .ZN(n248) );
  OA21D0 U241 ( .A1(N37), .A2(n256), .B(n242), .Z(n255) );
  CKND2D0 U242 ( .A1(N37), .A2(n256), .ZN(n242) );
  CKXOR2D0 U243 ( .A1(n241), .A2(n240), .Z(n256) );
  XNR2D0 U244 ( .A1(n257), .A2(n258), .ZN(n240) );
  NR2D0 U245 ( .A1(n259), .A2(n260), .ZN(n257) );
  XNR2D0 U246 ( .A1(n261), .A2(n262), .ZN(n241) );
  CKND2D0 U247 ( .A1(n263), .A2(n264), .ZN(n262) );
  OA21D0 U248 ( .A1(n265), .A2(n266), .B(n249), .Z(n254) );
  CKND2D0 U249 ( .A1(n265), .A2(n266), .ZN(n249) );
  OAI21D0 U250 ( .A1(n267), .A2(n268), .B(n269), .ZN(n266) );
  OA21D0 U251 ( .A1(n270), .A2(n271), .B(n247), .Z(n265) );
  CKND2D0 U252 ( .A1(n270), .A2(n271), .ZN(n247) );
  XNR2D0 U253 ( .A1(n272), .A2(n273), .ZN(n271) );
  CKND2D0 U254 ( .A1(n274), .A2(n275), .ZN(n273) );
  CKXOR2D0 U255 ( .A1(n245), .A2(n246), .Z(n270) );
  CKND2D0 U256 ( .A1(mantissa_b[9]), .A2(mantissa_a[1]), .ZN(n246) );
  XNR2D0 U257 ( .A1(n276), .A2(n277), .ZN(n245) );
  AN2D0 U258 ( .A1(n278), .A2(n279), .Z(n276) );
  XNR2D0 U259 ( .A1(n250), .A2(n251), .ZN(n252) );
  OA21D0 U260 ( .A1(n280), .A2(n281), .B(n282), .Z(n251) );
  AN2D0 U261 ( .A1(n283), .A2(n284), .Z(n250) );
  OAI21D0 U262 ( .A1(n285), .A2(n286), .B(n287), .ZN(N337) );
  CKXOR2D0 U263 ( .A1(n286), .A2(n285), .Z(N336) );
  OAI21D0 U264 ( .A1(n288), .A2(n289), .B(n283), .ZN(n285) );
  CKND2D0 U265 ( .A1(n288), .A2(n289), .ZN(n283) );
  OA21D0 U266 ( .A1(n290), .A2(n291), .B(n269), .Z(n289) );
  CKND2D0 U267 ( .A1(n290), .A2(n291), .ZN(n269) );
  CKXOR2D0 U268 ( .A1(n268), .A2(n267), .Z(n291) );
  XNR2D0 U269 ( .A1(n260), .A2(n259), .ZN(n267) );
  XNR2D0 U270 ( .A1(n263), .A2(n264), .ZN(n268) );
  CKXOR2D0 U271 ( .A1(n292), .A2(n293), .Z(n290) );
  OA21D0 U272 ( .A1(n294), .A2(n295), .B(n284), .Z(n288) );
  CKND2D0 U273 ( .A1(n294), .A2(n295), .ZN(n284) );
  OAI21D0 U274 ( .A1(n296), .A2(n297), .B(n298), .ZN(n295) );
  OA21D0 U275 ( .A1(n299), .A2(n300), .B(n282), .Z(n294) );
  CKND2D0 U276 ( .A1(n299), .A2(n300), .ZN(n282) );
  CKXOR2D0 U277 ( .A1(n280), .A2(n281), .Z(n300) );
  CKND2D0 U278 ( .A1(mantissa_b[9]), .A2(mantissa_a[0]), .ZN(n281) );
  CKXOR2D0 U279 ( .A1(n301), .A2(n278), .Z(n280) );
  CKXOR2D0 U280 ( .A1(n274), .A2(n275), .Z(n299) );
  OAI21D0 U281 ( .A1(n302), .A2(n303), .B(n287), .ZN(n286) );
  IND3D0 U282 ( .A1(n304), .B1(n305), .B2(n303), .ZN(n287) );
  CKND2D0 U283 ( .A1(n306), .A2(n307), .ZN(n303) );
  INR2D0 U284 ( .A1(n305), .B1(n304), .ZN(n302) );
  OAI21D0 U285 ( .A1(n308), .A2(n309), .B(n310), .ZN(N333) );
  CKND0 U286 ( .I(n38), .ZN(N332) );
  XNR2D0 U287 ( .A1(n309), .A2(n308), .ZN(n38) );
  OAI21D0 U288 ( .A1(n311), .A2(n312), .B(n306), .ZN(n308) );
  CKND2D0 U289 ( .A1(n311), .A2(n312), .ZN(n306) );
  OA21D0 U290 ( .A1(n313), .A2(n314), .B(n298), .Z(n312) );
  CKND2D0 U291 ( .A1(n313), .A2(n314), .ZN(n298) );
  CKXOR2D0 U292 ( .A1(n297), .A2(n296), .Z(n314) );
  CKXOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n296) );
  CKND2D0 U294 ( .A1(n317), .A2(n318), .ZN(n316) );
  XNR2D0 U295 ( .A1(n319), .A2(n320), .ZN(n297) );
  AN2D0 U296 ( .A1(n321), .A2(n322), .Z(n319) );
  XNR2D0 U297 ( .A1(n323), .A2(n324), .ZN(n313) );
  CKND2D0 U298 ( .A1(n325), .A2(n326), .ZN(n324) );
  OA21D0 U299 ( .A1(n327), .A2(n328), .B(n307), .Z(n311) );
  CKND2D0 U300 ( .A1(n327), .A2(n328), .ZN(n307) );
  OAI21D0 U301 ( .A1(n329), .A2(n330), .B(n331), .ZN(n328) );
  XNR2D0 U302 ( .A1(n304), .A2(n305), .ZN(n327) );
  CKXOR2D0 U303 ( .A1(n332), .A2(n333), .Z(n305) );
  INR2D0 U304 ( .A1(n334), .B1(n68), .ZN(n332) );
  XNR2D0 U305 ( .A1(n335), .A2(n336), .ZN(n304) );
  NR2D0 U306 ( .A1(n337), .A2(n338), .ZN(n335) );
  OAI21D0 U307 ( .A1(n339), .A2(n340), .B(n310), .ZN(n309) );
  IND3D0 U308 ( .A1(n341), .B1(n340), .B2(n342), .ZN(n310) );
  OAI21D0 U309 ( .A1(n343), .A2(n344), .B(n345), .ZN(n340) );
  INR2D0 U310 ( .A1(n342), .B1(n341), .ZN(n339) );
  CKND0 U311 ( .I(n42), .ZN(N329) );
  CKND2D0 U312 ( .A1(n346), .A2(n347), .ZN(n42) );
  CKXOR2D0 U313 ( .A1(n346), .A2(n347), .Z(N328) );
  OAI22D0 U314 ( .A1(n348), .A2(n349), .B1(n350), .B2(n351), .ZN(n347) );
  CKXOR2D0 U315 ( .A1(n344), .A2(n343), .Z(n346) );
  OAI21D0 U316 ( .A1(n352), .A2(n353), .B(n331), .ZN(n343) );
  CKND2D0 U317 ( .A1(n352), .A2(n353), .ZN(n331) );
  CKXOR2D0 U318 ( .A1(n330), .A2(n329), .Z(n353) );
  XNR2D0 U319 ( .A1(n317), .A2(n318), .ZN(n329) );
  CKXOR2D0 U320 ( .A1(n354), .A2(n321), .Z(n330) );
  CKXOR2D0 U321 ( .A1(n325), .A2(n326), .Z(n352) );
  OAI21D0 U322 ( .A1(n355), .A2(n356), .B(n345), .ZN(n344) );
  CKND2D0 U323 ( .A1(n355), .A2(n356), .ZN(n345) );
  OAI21D0 U324 ( .A1(n357), .A2(n358), .B(n359), .ZN(n356) );
  XNR2D0 U325 ( .A1(n342), .A2(n341), .ZN(n355) );
  CKXOR2D0 U326 ( .A1(n334), .A2(n68), .Z(n341) );
  CKXOR2D0 U327 ( .A1(n338), .A2(n337), .Z(n342) );
  CKND0 U328 ( .I(n41), .ZN(N327) );
  CKND2D0 U329 ( .A1(n360), .A2(n361), .ZN(n41) );
  CKXOR2D0 U330 ( .A1(n360), .A2(n361), .Z(N326) );
  OAI22D0 U331 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .ZN(n361) );
  CKXOR2D0 U332 ( .A1(n350), .A2(n351), .Z(n360) );
  OAI21D0 U333 ( .A1(n366), .A2(n367), .B(n359), .ZN(n351) );
  CKND2D0 U334 ( .A1(n366), .A2(n367), .ZN(n359) );
  CKXOR2D0 U335 ( .A1(n358), .A2(n357), .Z(n367) );
  XNR2D0 U336 ( .A1(n368), .A2(n369), .ZN(n357) );
  NR2D0 U337 ( .A1(n370), .A2(n371), .ZN(n368) );
  XNR2D0 U338 ( .A1(n372), .A2(n373), .ZN(n358) );
  CKND2D0 U339 ( .A1(n374), .A2(n375), .ZN(n373) );
  CKXOR2D0 U340 ( .A1(n376), .A2(n377), .Z(n366) );
  NR2D0 U341 ( .A1(n378), .A2(n379), .ZN(n376) );
  XNR2D0 U342 ( .A1(n348), .A2(n349), .ZN(n350) );
  XNR2D0 U343 ( .A1(n380), .A2(n381), .ZN(n349) );
  INR2D0 U344 ( .A1(n382), .B1(n73), .ZN(n380) );
  OA21D0 U345 ( .A1(n383), .A2(n384), .B(n385), .Z(n348) );
  INR3D0 U346 ( .A1(n386), .B1(n387), .B2(n388), .ZN(N325) );
  CKXOR2D0 U347 ( .A1(n388), .A2(n389), .Z(N324) );
  IND2D0 U348 ( .A1(n387), .B1(n386), .ZN(n389) );
  XNR2D0 U349 ( .A1(n364), .A2(n365), .ZN(n388) );
  OAI21D0 U350 ( .A1(n390), .A2(n391), .B(n385), .ZN(n365) );
  CKND2D0 U351 ( .A1(n390), .A2(n391), .ZN(n385) );
  CKXOR2D0 U352 ( .A1(n384), .A2(n383), .Z(n391) );
  XNR2D0 U353 ( .A1(n371), .A2(n370), .ZN(n383) );
  XNR2D0 U354 ( .A1(n374), .A2(n375), .ZN(n384) );
  CKXOR2D0 U355 ( .A1(n379), .A2(n378), .Z(n390) );
  XNR2D0 U356 ( .A1(n362), .A2(n363), .ZN(n364) );
  CKXOR2D0 U357 ( .A1(n382), .A2(n73), .Z(n363) );
  MAOI22D0 U358 ( .A1(n392), .A2(n393), .B1(n394), .B2(n395), .ZN(n362) );
  INR2D0 U359 ( .A1(n115), .B1(n116), .ZN(N323) );
  ND3D0 U360 ( .A1(n111), .A2(n108), .A3(n110), .ZN(n116) );
  CKXOR2D0 U361 ( .A1(n396), .A2(n397), .Z(n110) );
  NR2D0 U362 ( .A1(n114), .A2(n113), .ZN(n396) );
  CKXOR2D0 U363 ( .A1(n398), .A2(n399), .Z(n108) );
  CKXOR2D0 U364 ( .A1(n400), .A2(n401), .Z(n111) );
  NR2D0 U365 ( .A1(n112), .A2(n89), .ZN(n400) );
  XNR2D0 U366 ( .A1(n387), .A2(n386), .ZN(n115) );
  OAI22D0 U367 ( .A1(n402), .A2(n403), .B1(n399), .B2(n398), .ZN(n386) );
  XNR2D0 U368 ( .A1(n403), .A2(n402), .ZN(n398) );
  XNR2D0 U369 ( .A1(n404), .A2(n405), .ZN(n399) );
  XNR2D0 U370 ( .A1(n406), .A2(n407), .ZN(n403) );
  CKXOR2D0 U371 ( .A1(n408), .A2(n79), .Z(n402) );
  XNR2D0 U372 ( .A1(n392), .A2(n393), .ZN(n387) );
  CKXOR2D0 U373 ( .A1(n409), .A2(n410), .Z(n393) );
  CKND2D0 U374 ( .A1(n404), .A2(n405), .ZN(n410) );
  CKXOR2D0 U375 ( .A1(n395), .A2(n394), .Z(n392) );
  XNR2D0 U376 ( .A1(n411), .A2(n412), .ZN(n394) );
  INR2D0 U377 ( .A1(n408), .B1(n79), .ZN(n411) );
  XNR2D0 U378 ( .A1(n413), .A2(n414), .ZN(n395) );
  NR2D0 U379 ( .A1(n407), .A2(n406), .ZN(n413) );
  OAI22D0 U380 ( .A1(n415), .A2(n416), .B1(n119), .B2(n120), .ZN(N317) );
  OAI21D0 U381 ( .A1(N37), .A2(n156), .B(n157), .ZN(n120) );
  CKXOR2D0 U382 ( .A1(N251), .A2(n416), .Z(n119) );
  CKXOR2D0 U383 ( .A1(n417), .A2(N118), .Z(n416) );
  CKND0 U384 ( .I(N251), .ZN(n415) );
  OAI21D0 U385 ( .A1(n418), .A2(n417), .B(n419), .ZN(N255) );
  OAI21D0 U386 ( .A1(n420), .A2(n421), .B(n419), .ZN(n417) );
  ND3D0 U387 ( .A1(mantissa_a[8]), .A2(n421), .A3(mantissa_b[9]), .ZN(n419) );
  CKXOR2D0 U388 ( .A1(n422), .A2(n423), .Z(n421) );
  NR2D0 U389 ( .A1(n70), .A2(n68), .ZN(n420) );
  CKND0 U390 ( .I(mantissa_a[8]), .ZN(n70) );
  OAI21D0 U391 ( .A1(n107), .A2(n106), .B(n157), .ZN(N251) );
  CKND2D0 U392 ( .A1(n156), .A2(N37), .ZN(n157) );
  IAO21D0 U393 ( .A1(n293), .A2(n292), .B(n99), .ZN(N37) );
  ND3D0 U394 ( .A1(n326), .A2(n325), .A3(n323), .ZN(n292) );
  XNR2D0 U395 ( .A1(n424), .A2(mantissa_b[1]), .ZN(n323) );
  AOI22D0 U396 ( .A1(mantissa_a[8]), .A2(n425), .B1(mantissa_a[9]), .B2(
        mantissa_b[0]), .ZN(n424) );
  INR3D0 U397 ( .A1(n377), .B1(n378), .B2(n379), .ZN(n325) );
  IND3D0 U398 ( .A1(n409), .B1(n405), .B2(n404), .ZN(n379) );
  INR3D0 U399 ( .A1(n397), .B1(n114), .B2(n113), .ZN(n404) );
  IND2D0 U400 ( .A1(n101), .B1(n100), .ZN(n113) );
  INR2D0 U401 ( .A1(n105), .B1(n99), .ZN(n100) );
  IND2D0 U402 ( .A1(n425), .B1(n426), .ZN(n105) );
  MUX2ND0 U403 ( .I0(n427), .I1(n102), .S(mantissa_b[1]), .ZN(n426) );
  NR2D0 U404 ( .A1(n102), .A2(n104), .ZN(n427) );
  CKND0 U405 ( .I(mantissa_b[0]), .ZN(n104) );
  CKND0 U406 ( .I(mantissa_a[0]), .ZN(n102) );
  XNR2D0 U407 ( .A1(n428), .A2(n99), .ZN(n101) );
  AOI22D0 U408 ( .A1(n425), .A2(mantissa_a[0]), .B1(mantissa_b[0]), .B2(
        mantissa_a[1]), .ZN(n428) );
  CKXOR2D0 U409 ( .A1(n429), .A2(mantissa_b[1]), .Z(n114) );
  AOI22D0 U410 ( .A1(n425), .A2(mantissa_a[1]), .B1(mantissa_b[0]), .B2(
        mantissa_a[2]), .ZN(n429) );
  CKXOR2D0 U411 ( .A1(n430), .A2(n99), .Z(n397) );
  AOI22D0 U412 ( .A1(n425), .A2(mantissa_a[2]), .B1(mantissa_b[0]), .B2(
        mantissa_a[3]), .ZN(n430) );
  CKXOR2D0 U413 ( .A1(n431), .A2(n99), .Z(n405) );
  AOI22D0 U414 ( .A1(n425), .A2(mantissa_a[3]), .B1(mantissa_b[0]), .B2(
        mantissa_a[4]), .ZN(n431) );
  XNR2D0 U415 ( .A1(n432), .A2(n99), .ZN(n409) );
  AOI22D0 U416 ( .A1(n425), .A2(mantissa_a[4]), .B1(mantissa_b[0]), .B2(
        mantissa_a[5]), .ZN(n432) );
  CKXOR2D0 U417 ( .A1(n433), .A2(mantissa_b[1]), .Z(n378) );
  AOI22D0 U418 ( .A1(n425), .A2(mantissa_a[5]), .B1(mantissa_b[0]), .B2(
        mantissa_a[6]), .ZN(n433) );
  CKXOR2D0 U455 ( .A1(n434), .A2(n99), .Z(n377) );
  AOI22D0 U456 ( .A1(n425), .A2(mantissa_a[6]), .B1(mantissa_a[7]), .B2(
        mantissa_b[0]), .ZN(n434) );
  CKXOR2D0 U457 ( .A1(n435), .A2(n99), .Z(n326) );
  AOI22D0 U458 ( .A1(mantissa_a[7]), .A2(n425), .B1(mantissa_a[8]), .B2(
        mantissa_b[0]), .ZN(n435) );
  NR2D0 U459 ( .A1(n99), .A2(mantissa_b[0]), .ZN(n425) );
  OAI21D0 U460 ( .A1(mantissa_b[0]), .A2(n66), .B(mantissa_b[1]), .ZN(n293) );
  CKXOR2D0 U461 ( .A1(n107), .A2(n106), .Z(n156) );
  OAI21D0 U462 ( .A1(n185), .A2(n184), .B(mantissa_b[5]), .ZN(n106) );
  ND3D0 U463 ( .A1(n208), .A2(n207), .A3(n205), .ZN(n184) );
  XNR2D0 U464 ( .A1(n436), .A2(mantissa_b[5]), .ZN(n205) );
  AOI22D0 U465 ( .A1(mantissa_a[9]), .A2(n437), .B1(mantissa_a[8]), .B2(n438), 
        .ZN(n436) );
  INR3D0 U466 ( .A1(n258), .B1(n259), .B2(n260), .ZN(n207) );
  ND3D0 U467 ( .A1(n318), .A2(n317), .A3(n315), .ZN(n260) );
  XNR2D0 U468 ( .A1(n439), .A2(mantissa_b[5]), .ZN(n315) );
  AOI22D0 U469 ( .A1(mantissa_a[5]), .A2(n437), .B1(n438), .B2(mantissa_a[4]), 
        .ZN(n439) );
  INR3D0 U470 ( .A1(n369), .B1(n370), .B2(n371), .ZN(n317) );
  ND3D0 U471 ( .A1(mantissa_b[5]), .A2(n408), .A3(n412), .ZN(n371) );
  CKXOR2D0 U472 ( .A1(n440), .A2(n79), .Z(n412) );
  AOI22D0 U473 ( .A1(mantissa_a[1]), .A2(n437), .B1(n438), .B2(mantissa_a[0]), 
        .ZN(n440) );
  XNR2D0 U474 ( .A1(mantissa_b[5]), .A2(n441), .ZN(n408) );
  CKND2D0 U475 ( .A1(mantissa_a[0]), .A2(n437), .ZN(n441) );
  XNR2D0 U476 ( .A1(n442), .A2(n79), .ZN(n370) );
  AOI22D0 U477 ( .A1(mantissa_a[2]), .A2(n437), .B1(n438), .B2(mantissa_a[1]), 
        .ZN(n442) );
  CKXOR2D0 U478 ( .A1(n443), .A2(n79), .Z(n369) );
  AOI22D0 U479 ( .A1(mantissa_a[3]), .A2(n437), .B1(n438), .B2(mantissa_a[2]), 
        .ZN(n443) );
  CKXOR2D0 U480 ( .A1(n444), .A2(n79), .Z(n318) );
  AOI22D0 U481 ( .A1(mantissa_a[4]), .A2(n437), .B1(n438), .B2(mantissa_a[3]), 
        .ZN(n444) );
  XNR2D0 U482 ( .A1(n445), .A2(n79), .ZN(n259) );
  AOI22D0 U483 ( .A1(mantissa_a[6]), .A2(n437), .B1(n438), .B2(mantissa_a[5]), 
        .ZN(n445) );
  CKXOR2D0 U484 ( .A1(n446), .A2(n79), .Z(n258) );
  AOI22D0 U485 ( .A1(mantissa_a[7]), .A2(n437), .B1(n438), .B2(mantissa_a[6]), 
        .ZN(n446) );
  CKXOR2D0 U486 ( .A1(n447), .A2(n79), .Z(n208) );
  AOI22D0 U487 ( .A1(mantissa_a[8]), .A2(n437), .B1(mantissa_a[7]), .B2(n438), 
        .ZN(n447) );
  CKXOR2D0 U488 ( .A1(n89), .A2(n84), .Z(n437) );
  CKND0 U489 ( .I(mantissa_b[4]), .ZN(n84) );
  CKXOR2D0 U490 ( .A1(mantissa_b[5]), .A2(n448), .Z(n185) );
  CKND2D0 U491 ( .A1(mantissa_a[9]), .A2(n438), .ZN(n448) );
  OA21D0 U492 ( .A1(mantissa_b[4]), .A2(n89), .B(n449), .Z(n438) );
  MUX2ND0 U493 ( .I0(n89), .I1(mantissa_b[4]), .S(mantissa_b[5]), .ZN(n449) );
  OAI21D0 U494 ( .A1(n237), .A2(n236), .B(mantissa_b[3]), .ZN(n107) );
  IND3D0 U495 ( .A1(n261), .B1(n264), .B2(n263), .ZN(n236) );
  AN3D0 U496 ( .A1(n322), .A2(n321), .A3(n320), .Z(n263) );
  CKXOR2D0 U497 ( .A1(n450), .A2(n89), .Z(n320) );
  AOI22D0 U498 ( .A1(mantissa_a[7]), .A2(n451), .B1(mantissa_a[6]), .B2(n452), 
        .ZN(n450) );
  CKXOR2D0 U499 ( .A1(n453), .A2(n89), .Z(n321) );
  AOI22D0 U500 ( .A1(mantissa_a[6]), .A2(n451), .B1(mantissa_a[5]), .B2(n452), 
        .ZN(n453) );
  CKND0 U501 ( .I(n354), .ZN(n322) );
  IND3D0 U502 ( .A1(n372), .B1(n375), .B2(n374), .ZN(n354) );
  INR3D0 U503 ( .A1(n414), .B1(n407), .B2(n406), .ZN(n374) );
  IND3D0 U504 ( .A1(n112), .B1(n401), .B2(mantissa_b[3]), .ZN(n406) );
  CKXOR2D0 U505 ( .A1(n454), .A2(n89), .Z(n401) );
  AOI22D0 U506 ( .A1(mantissa_a[1]), .A2(n451), .B1(n452), .B2(mantissa_a[0]), 
        .ZN(n454) );
  CKXOR2D0 U507 ( .A1(mantissa_b[3]), .A2(n455), .Z(n112) );
  CKND2D0 U508 ( .A1(mantissa_a[0]), .A2(n451), .ZN(n455) );
  XNR2D0 U509 ( .A1(n456), .A2(n89), .ZN(n407) );
  AOI22D0 U510 ( .A1(mantissa_a[2]), .A2(n451), .B1(n452), .B2(mantissa_a[1]), 
        .ZN(n456) );
  CKXOR2D0 U511 ( .A1(n457), .A2(n89), .Z(n414) );
  AOI22D0 U512 ( .A1(mantissa_a[3]), .A2(n451), .B1(mantissa_a[2]), .B2(n452), 
        .ZN(n457) );
  CKXOR2D0 U513 ( .A1(n458), .A2(n89), .Z(n375) );
  AOI22D0 U514 ( .A1(mantissa_a[4]), .A2(n451), .B1(mantissa_a[3]), .B2(n452), 
        .ZN(n458) );
  XNR2D0 U515 ( .A1(n459), .A2(n89), .ZN(n372) );
  AOI22D0 U516 ( .A1(mantissa_a[5]), .A2(n451), .B1(mantissa_a[4]), .B2(n452), 
        .ZN(n459) );
  CKXOR2D0 U517 ( .A1(n460), .A2(n89), .Z(n264) );
  AOI22D0 U518 ( .A1(mantissa_a[8]), .A2(n451), .B1(mantissa_a[7]), .B2(n452), 
        .ZN(n460) );
  XNR2D0 U519 ( .A1(n461), .A2(n89), .ZN(n261) );
  CKND0 U520 ( .I(mantissa_b[3]), .ZN(n89) );
  AOI22D0 U521 ( .A1(mantissa_a[9]), .A2(n451), .B1(mantissa_a[8]), .B2(n452), 
        .ZN(n461) );
  CKXOR2D0 U522 ( .A1(n99), .A2(n94), .Z(n451) );
  CKND0 U523 ( .I(mantissa_b[2]), .ZN(n94) );
  CKXOR2D0 U524 ( .A1(mantissa_b[3]), .A2(n462), .Z(n237) );
  CKND2D0 U525 ( .A1(mantissa_a[9]), .A2(n452), .ZN(n462) );
  OA21D0 U526 ( .A1(mantissa_b[2]), .A2(n99), .B(n463), .Z(n452) );
  MUX2ND0 U527 ( .I0(n99), .I1(mantissa_b[2]), .S(mantissa_b[3]), .ZN(n463) );
  CKND0 U528 ( .I(mantissa_b[1]), .ZN(n99) );
  NR2D0 U529 ( .A1(n68), .A2(n66), .ZN(N142) );
  AOI21D0 U530 ( .A1(n422), .A2(n423), .B(n68), .ZN(N141) );
  XNR2D0 U531 ( .A1(n464), .A2(n68), .ZN(n423) );
  NR2D0 U532 ( .A1(n465), .A2(n66), .ZN(n464) );
  CKND0 U533 ( .I(mantissa_a[9]), .ZN(n66) );
  AN3D0 U534 ( .A1(n132), .A2(n135), .A3(n134), .Z(n422) );
  AN3D0 U535 ( .A1(n170), .A2(n171), .A3(n169), .Z(n134) );
  CKXOR2D0 U536 ( .A1(n466), .A2(n68), .Z(n169) );
  AOI22D0 U537 ( .A1(mantissa_a[6]), .A2(n467), .B1(mantissa_a[7]), .B2(n468), 
        .ZN(n466) );
  CKND0 U538 ( .I(n192), .ZN(n171) );
  IND3D0 U539 ( .A1(n220), .B1(n223), .B2(n222), .ZN(n192) );
  AN3D0 U540 ( .A1(n278), .A2(n279), .A3(n277), .Z(n222) );
  CKXOR2D0 U541 ( .A1(n469), .A2(n68), .Z(n277) );
  AOI22D0 U542 ( .A1(mantissa_a[2]), .A2(n467), .B1(mantissa_a[3]), .B2(n468), 
        .ZN(n469) );
  CKND0 U543 ( .I(n301), .ZN(n279) );
  ND3D0 U544 ( .A1(mantissa_b[9]), .A2(n334), .A3(n333), .ZN(n301) );
  CKXOR2D0 U545 ( .A1(n470), .A2(n68), .Z(n333) );
  AOI22D0 U546 ( .A1(mantissa_a[0]), .A2(n467), .B1(mantissa_a[1]), .B2(n468), 
        .ZN(n470) );
  XNR2D0 U547 ( .A1(mantissa_b[9]), .A2(n471), .ZN(n334) );
  CKND2D0 U548 ( .A1(mantissa_a[0]), .A2(n468), .ZN(n471) );
  CKXOR2D0 U549 ( .A1(n472), .A2(n68), .Z(n278) );
  AOI22D0 U550 ( .A1(mantissa_a[1]), .A2(n467), .B1(mantissa_a[2]), .B2(n468), 
        .ZN(n472) );
  CKXOR2D0 U551 ( .A1(n473), .A2(n68), .Z(n223) );
  AOI22D0 U552 ( .A1(mantissa_a[3]), .A2(n467), .B1(mantissa_a[4]), .B2(n468), 
        .ZN(n473) );
  XNR2D0 U553 ( .A1(n474), .A2(n68), .ZN(n220) );
  AOI22D0 U554 ( .A1(mantissa_a[4]), .A2(n467), .B1(mantissa_a[5]), .B2(n468), 
        .ZN(n474) );
  CKXOR2D0 U555 ( .A1(n475), .A2(n68), .Z(n170) );
  AOI22D0 U556 ( .A1(mantissa_a[5]), .A2(n467), .B1(mantissa_a[6]), .B2(n468), 
        .ZN(n475) );
  CKXOR2D0 U557 ( .A1(n476), .A2(n68), .Z(n135) );
  CKND0 U558 ( .I(mantissa_b[9]), .ZN(n68) );
  AOI22D0 U559 ( .A1(mantissa_a[7]), .A2(n467), .B1(mantissa_a[8]), .B2(n468), 
        .ZN(n476) );
  XNR2D0 U560 ( .A1(n477), .A2(mantissa_b[9]), .ZN(n132) );
  AOI22D0 U561 ( .A1(mantissa_a[8]), .A2(n467), .B1(mantissa_a[9]), .B2(n468), 
        .ZN(n477) );
  CKXOR2D0 U562 ( .A1(n73), .A2(n71), .Z(n468) );
  CKND0 U563 ( .I(n465), .ZN(n467) );
  MUX2ND0 U564 ( .I0(n478), .I1(n479), .S(mantissa_b[9]), .ZN(n465) );
  NR2D0 U565 ( .A1(mantissa_b[8]), .A2(mantissa_b[7]), .ZN(n479) );
  NR2D0 U566 ( .A1(n73), .A2(n71), .ZN(n478) );
  CKND0 U567 ( .I(mantissa_b[8]), .ZN(n71) );
  CKND0 U568 ( .I(n418), .ZN(N118) );
  OAI21D0 U569 ( .A1(n130), .A2(n131), .B(mantissa_b[7]), .ZN(n418) );
  ND3D0 U570 ( .A1(n167), .A2(n166), .A3(n164), .ZN(n131) );
  XNR2D0 U571 ( .A1(n480), .A2(mantissa_b[7]), .ZN(n164) );
  AOI22D0 U572 ( .A1(mantissa_a[9]), .A2(n481), .B1(n482), .B2(mantissa_a[8]), 
        .ZN(n480) );
  INR3D0 U573 ( .A1(n217), .B1(n218), .B2(n219), .ZN(n166) );
  ND3D0 U574 ( .A1(n275), .A2(n274), .A3(n272), .ZN(n219) );
  XNR2D0 U575 ( .A1(n483), .A2(mantissa_b[7]), .ZN(n272) );
  AOI22D0 U576 ( .A1(mantissa_a[5]), .A2(n481), .B1(n482), .B2(mantissa_a[4]), 
        .ZN(n483) );
  INR3D0 U577 ( .A1(n336), .B1(n337), .B2(n338), .ZN(n274) );
  ND3D0 U578 ( .A1(mantissa_b[7]), .A2(n382), .A3(n381), .ZN(n338) );
  CKXOR2D0 U579 ( .A1(n484), .A2(n73), .Z(n381) );
  AOI22D0 U580 ( .A1(mantissa_a[1]), .A2(n481), .B1(n482), .B2(mantissa_a[0]), 
        .ZN(n484) );
  XNR2D0 U581 ( .A1(mantissa_b[7]), .A2(n485), .ZN(n382) );
  CKND2D0 U582 ( .A1(mantissa_a[0]), .A2(n481), .ZN(n485) );
  XNR2D0 U583 ( .A1(n486), .A2(n73), .ZN(n337) );
  AOI22D0 U584 ( .A1(mantissa_a[2]), .A2(n481), .B1(n482), .B2(mantissa_a[1]), 
        .ZN(n486) );
  CKXOR2D0 U585 ( .A1(n487), .A2(n73), .Z(n336) );
  AOI22D0 U586 ( .A1(mantissa_a[3]), .A2(n481), .B1(n482), .B2(mantissa_a[2]), 
        .ZN(n487) );
  CKXOR2D0 U587 ( .A1(n488), .A2(n73), .Z(n275) );
  AOI22D0 U588 ( .A1(mantissa_a[4]), .A2(n481), .B1(n482), .B2(mantissa_a[3]), 
        .ZN(n488) );
  CKXOR2D0 U589 ( .A1(n489), .A2(mantissa_b[7]), .Z(n218) );
  AOI22D0 U590 ( .A1(mantissa_a[6]), .A2(n481), .B1(n482), .B2(mantissa_a[5]), 
        .ZN(n489) );
  CKXOR2D0 U591 ( .A1(n490), .A2(n73), .Z(n217) );
  AOI22D0 U592 ( .A1(mantissa_a[7]), .A2(n481), .B1(n482), .B2(mantissa_a[6]), 
        .ZN(n490) );
  CKXOR2D0 U593 ( .A1(n491), .A2(n73), .Z(n167) );
  CKND0 U594 ( .I(mantissa_b[7]), .ZN(n73) );
  AOI22D0 U595 ( .A1(mantissa_a[8]), .A2(n481), .B1(n482), .B2(mantissa_a[7]), 
        .ZN(n491) );
  XNR2D0 U596 ( .A1(n79), .A2(mantissa_b[6]), .ZN(n481) );
  CKXOR2D0 U597 ( .A1(mantissa_b[7]), .A2(n492), .Z(n130) );
  CKND2D0 U598 ( .A1(mantissa_a[9]), .A2(n482), .ZN(n492) );
  OA21D0 U599 ( .A1(mantissa_b[6]), .A2(n79), .B(n493), .Z(n482) );
  MUX2ND0 U600 ( .I0(n79), .I1(mantissa_b[6]), .S(mantissa_b[7]), .ZN(n493) );
  CKND0 U601 ( .I(mantissa_b[5]), .ZN(n79) );
endmodule


module fma_lza_1 ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, 
        sign_ab, sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  assign lza_done = adder_start;

  NR2D0 U3 ( .A1(n168), .A2(n169), .ZN(mantissa_shift[4]) );
  CKXOR2D0 U4 ( .A1(n170), .A2(n171), .Z(n169) );
  NR2D0 U5 ( .A1(n172), .A2(n173), .ZN(n170) );
  AOI21D0 U6 ( .A1(n174), .A2(n175), .B(n168), .ZN(mantissa_shift[3]) );
  IND2D0 U7 ( .A1(n173), .B1(n176), .ZN(n175) );
  MUX2ND0 U8 ( .I0(n177), .I1(n172), .S(n173), .ZN(n174) );
  OAI21D0 U9 ( .A1(n178), .A2(n179), .B(n180), .ZN(n173) );
  NR2D0 U10 ( .A1(n176), .A2(n177), .ZN(n172) );
  AN2D0 U11 ( .A1(n181), .A2(n182), .Z(n176) );
  MUX2ND0 U12 ( .I0(n183), .I1(n184), .S(n185), .ZN(n181) );
  AOI221D0 U13 ( .A1(n186), .A2(n187), .B1(n188), .B2(n189), .C(n171), .ZN(
        n177) );
  MUX2D0 U14 ( .I0(n190), .I1(n191), .S(sign_c), .Z(n171) );
  NR2D0 U15 ( .A1(n186), .A2(n187), .ZN(n191) );
  NR2D0 U16 ( .A1(n188), .A2(n189), .ZN(n190) );
  IOA21D0 U17 ( .A1(n192), .A2(n193), .B(n194), .ZN(n189) );
  OAI21D0 U18 ( .A1(n195), .A2(n186), .B(n196), .ZN(n187) );
  NR2D0 U19 ( .A1(n168), .A2(n197), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U20 ( .A1(n198), .A2(n178), .Z(n197) );
  MUX2D0 U21 ( .I0(n199), .I1(n200), .S(sign_c), .Z(n178) );
  CKXOR2D0 U22 ( .A1(n201), .A2(n202), .Z(n200) );
  AOI21D0 U23 ( .A1(n203), .A2(n204), .B(n183), .ZN(n201) );
  CKND2D0 U24 ( .A1(n205), .A2(n206), .ZN(n183) );
  XNR2D0 U25 ( .A1(n207), .A2(n208), .ZN(n199) );
  IND2D0 U26 ( .A1(n184), .B1(n209), .ZN(n208) );
  CKND2D0 U27 ( .A1(n210), .A2(n211), .ZN(n184) );
  NR2D0 U28 ( .A1(n179), .A2(n212), .ZN(n198) );
  MUX2D0 U29 ( .I0(n213), .I1(n214), .S(sign_c), .Z(n179) );
  CKXOR2D0 U30 ( .A1(n196), .A2(n215), .Z(n214) );
  OR2D0 U31 ( .A1(n186), .A2(n195), .Z(n215) );
  AOI21D0 U32 ( .A1(n216), .A2(n217), .B(n218), .ZN(n196) );
  CKXOR2D0 U33 ( .A1(n194), .A2(n219), .Z(n213) );
  CKND2D0 U34 ( .A1(n193), .A2(n192), .ZN(n219) );
  CKND2D0 U35 ( .A1(n220), .A2(n221), .ZN(n192) );
  AOI21D0 U36 ( .A1(n222), .A2(n223), .B(n224), .ZN(n194) );
  AOI211D0 U37 ( .A1(n212), .A2(n225), .B(n226), .C(n168), .ZN(
        mantissa_shift[1]) );
  MUX2ND0 U38 ( .I0(n227), .I1(n228), .S(n185), .ZN(n226) );
  CKND2D0 U39 ( .A1(n229), .A2(n222), .ZN(n228) );
  OAI21D0 U40 ( .A1(n230), .A2(n231), .B(n188), .ZN(n222) );
  CKND0 U41 ( .I(n193), .ZN(n188) );
  NR2D0 U42 ( .A1(n232), .A2(n233), .ZN(n193) );
  NR2D0 U43 ( .A1(n234), .A2(n232), .ZN(n230) );
  NR2D0 U44 ( .A1(n235), .A2(n236), .ZN(n232) );
  CKXOR2D0 U45 ( .A1(n223), .A2(n224), .Z(n229) );
  NR2D0 U46 ( .A1(n237), .A2(n235), .ZN(n224) );
  AN2D0 U47 ( .A1(n238), .A2(n239), .Z(n223) );
  CKND2D0 U48 ( .A1(n240), .A2(n216), .ZN(n227) );
  OAI21D0 U49 ( .A1(n241), .A2(n242), .B(n186), .ZN(n216) );
  CKND2D0 U50 ( .A1(n242), .A2(n241), .ZN(n186) );
  CKXOR2D0 U51 ( .A1(n217), .A2(n218), .Z(n240) );
  IAO21D0 U52 ( .A1(n243), .A2(n195), .B(n244), .ZN(n217) );
  INR2D0 U53 ( .A1(n245), .B1(n246), .ZN(n195) );
  INR2D0 U54 ( .A1(n246), .B1(n245), .ZN(n243) );
  ND3D0 U55 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  CKND0 U56 ( .I(n180), .ZN(n212) );
  AOI21D0 U57 ( .A1(n248), .A2(n247), .B(n249), .ZN(n180) );
  AN2D0 U58 ( .A1(n250), .A2(n182), .Z(n249) );
  MUX2D0 U59 ( .I0(n207), .I1(n202), .S(sign_c), .Z(n182) );
  CKND2D0 U60 ( .A1(n251), .A2(n252), .ZN(n202) );
  XNR2D0 U61 ( .A1(n205), .A2(n206), .ZN(n251) );
  CKND2D0 U62 ( .A1(n253), .A2(n254), .ZN(n207) );
  XNR2D0 U63 ( .A1(n211), .A2(n210), .ZN(n254) );
  MUX2ND0 U64 ( .I0(n255), .I1(n256), .S(n185), .ZN(n250) );
  CKND2D0 U65 ( .A1(n257), .A2(n258), .ZN(n256) );
  OAI21D0 U66 ( .A1(n259), .A2(n260), .B(n209), .ZN(n258) );
  CKND2D0 U67 ( .A1(n259), .A2(n260), .ZN(n209) );
  IND3D0 U68 ( .A1(n261), .B1(n262), .B2(n263), .ZN(n255) );
  XNR2D0 U69 ( .A1(n203), .A2(n204), .ZN(n262) );
  NR2D0 U70 ( .A1(n264), .A2(n168), .ZN(mantissa_shift[0]) );
  OR2D0 U71 ( .A1(fma_byp), .A2(sign_ab), .Z(n168) );
  XNR2D0 U72 ( .A1(n248), .A2(n247), .ZN(n264) );
  MUX2ND0 U73 ( .I0(n265), .I1(n266), .S(n185), .ZN(n247) );
  AOI22D0 U74 ( .A1(n259), .A2(n267), .B1(n210), .B2(n268), .ZN(n266) );
  OAI21D0 U75 ( .A1(n253), .A2(n269), .B(n270), .ZN(n268) );
  IAO21D0 U76 ( .A1(n271), .A2(n272), .B(n273), .ZN(n210) );
  OAI31D0 U77 ( .A1(n257), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B(n274), 
        .ZN(n267) );
  AOI21D0 U78 ( .A1(n260), .A2(n275), .B(n276), .ZN(n259) );
  AOI22D0 U79 ( .A1(n203), .A2(n277), .B1(n205), .B2(n278), .ZN(n265) );
  OAI21D0 U80 ( .A1(n279), .A2(n280), .B(n281), .ZN(n278) );
  CKND0 U81 ( .I(n282), .ZN(n279) );
  MUX2ND0 U82 ( .I0(n283), .I1(n284), .S(n206), .ZN(n205) );
  NR3D0 U83 ( .A1(n285), .A2(n281), .A3(n286), .ZN(n284) );
  OAI21D0 U84 ( .A1(n263), .A2(n261), .B(n287), .ZN(n277) );
  CKND0 U85 ( .I(n288), .ZN(n287) );
  CKND0 U86 ( .I(n289), .ZN(n263) );
  CKND2D0 U87 ( .A1(n290), .A2(n291), .ZN(n203) );
  OAI21D0 U88 ( .A1(n292), .A2(n293), .B(n294), .ZN(n291) );
  OAI31D0 U89 ( .A1(n185), .A2(n218), .A3(n295), .B(n296), .ZN(n248) );
  MUX2ND0 U90 ( .I0(n235), .I1(n297), .S(n236), .ZN(n296) );
  AOI21D0 U91 ( .A1(n231), .A2(n298), .B(n299), .ZN(n236) );
  CKXOR2D0 U92 ( .A1(n237), .A2(n235), .Z(n297) );
  CKND2D0 U93 ( .A1(n220), .A2(n300), .ZN(n237) );
  OAI21D0 U94 ( .A1(n238), .A2(n301), .B(n302), .ZN(n300) );
  XNR2D0 U95 ( .A1(n239), .A2(n221), .ZN(n220) );
  OR2D0 U96 ( .A1(n303), .A2(n304), .Z(n239) );
  ND4D0 U97 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n235) );
  NR4D0 U98 ( .A1(n309), .A2(n310), .A3(n234), .A4(n311), .ZN(n308) );
  OAI31D0 U99 ( .A1(n303), .A2(n312), .A3(n313), .B(n261), .ZN(n311) );
  INR3D0 U100 ( .A1(n299), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n234)
         );
  AO31D0 U101 ( .A1(n275), .A2(mantissa_ab[17]), .A3(mantissa_c[17]), .B(n314), 
        .Z(n310) );
  AO33D0 U102 ( .A1(mantissa_c[2]), .A2(mantissa_ab[2]), .A3(n298), .B1(
        mantissa_c[3]), .B2(mantissa_ab[3]), .B3(n304), .Z(n314) );
  OAI211D0 U103 ( .A1(n272), .A2(n315), .B(n316), .C(n317), .ZN(n309) );
  AOI31D0 U104 ( .A1(mantissa_c[8]), .A2(mantissa_ab[8]), .A3(n318), .B(n319), 
        .ZN(n317) );
  AO33D0 U105 ( .A1(n320), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B1(n253), .B2(mantissa_ab[13]), .B3(mantissa_c[13]), .Z(n319) );
  CKND0 U106 ( .I(n301), .ZN(n318) );
  AOI33D0 U107 ( .A1(mantissa_c[0]), .A2(mantissa_ab[0]), .A3(n299), .B1(
        mantissa_c[15]), .B2(mantissa_ab[15]), .B3(n276), .ZN(n316) );
  NR3D0 U108 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n231), .ZN(n299)
         );
  CKND0 U109 ( .I(n233), .ZN(n231) );
  CKND2D0 U110 ( .A1(mantissa_c[11]), .A2(mantissa_ab[11]), .ZN(n315) );
  AOI211D0 U111 ( .A1(n271), .A2(n283), .B(n321), .C(n322), .ZN(n307) );
  OAI33D0 U112 ( .A1(n289), .A2(mantissa_c[21]), .A3(mantissa_ab[21]), .B1(
        n270), .B2(n286), .B3(n285), .ZN(n322) );
  CKND0 U113 ( .I(n323), .ZN(n270) );
  OAI31D0 U114 ( .A1(n324), .A2(n325), .A3(n326), .B(n327), .ZN(n321) );
  AOI33D0 U115 ( .A1(mantissa_c[1]), .A2(mantissa_ab[1]), .A3(n233), .B1(
        mantissa_c[9]), .B2(mantissa_ab[9]), .B3(n273), .ZN(n327) );
  INR3D0 U116 ( .A1(n298), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n233)
         );
  INR3D0 U117 ( .A1(n304), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n298)
         );
  NR3D0 U118 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n221), .ZN(n304)
         );
  CKND0 U119 ( .I(n328), .ZN(n221) );
  AOI31D0 U120 ( .A1(mantissa_c[7]), .A2(mantissa_ab[7]), .A3(n238), .B(n329), 
        .ZN(n306) );
  OAI32D0 U121 ( .A1(n260), .A2(n292), .A3(n293), .B1(n282), .B2(n269), .ZN(
        n329) );
  CKND0 U122 ( .I(mantissa_ab[16]), .ZN(n292) );
  AOI33D0 U123 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n330), .B1(
        mantissa_c[4]), .B2(mantissa_ab[4]), .B3(n328), .ZN(n305) );
  NR3D0 U124 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n303), .ZN(n328)
         );
  OR3D0 U125 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n302), .Z(n303) );
  CKND0 U126 ( .I(n302), .ZN(n330) );
  ND3D0 U127 ( .A1(n331), .A2(n332), .A3(n238), .ZN(n302) );
  NR3D0 U128 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n301), .ZN(n238)
         );
  ND3D0 U129 ( .A1(n333), .A2(n334), .A3(n273), .ZN(n301) );
  NR3D0 U130 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n211), .ZN(n273)
         );
  CKND0 U131 ( .I(n271), .ZN(n211) );
  NR3D0 U132 ( .A1(mantissa_ab[11]), .A2(mantissa_c[11]), .A3(n272), .ZN(n271)
         );
  ND3D0 U133 ( .A1(n286), .A2(n285), .A3(n323), .ZN(n272) );
  INR3D0 U134 ( .A1(n253), .B1(mantissa_ab[13]), .B2(mantissa_c[13]), .ZN(n323) );
  NR3D0 U135 ( .A1(mantissa_ab[14]), .A2(mantissa_c[14]), .A3(n269), .ZN(n253)
         );
  IND3D0 U136 ( .A1(mantissa_ab[15]), .B1(n276), .B2(n335), .ZN(n269) );
  NR3D0 U137 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n260), .ZN(n276)
         );
  CKND0 U138 ( .I(n336), .ZN(n260) );
  INR3D0 U139 ( .A1(n275), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n336) );
  NR3D0 U140 ( .A1(mantissa_ab[18]), .A2(mantissa_c[18]), .A3(n274), .ZN(n275)
         );
  CKND0 U141 ( .I(n320), .ZN(n274) );
  NR3D0 U142 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n324), .ZN(n320)
         );
  CKND0 U143 ( .I(n257), .ZN(n324) );
  NR4D0 U144 ( .A1(mantissa_ab[20]), .A2(mantissa_ab[21]), .A3(mantissa_c[20]), 
        .A4(mantissa_c[21]), .ZN(n257) );
  CKND0 U145 ( .I(mantissa_c[12]), .ZN(n285) );
  CKND0 U146 ( .I(mantissa_ab[12]), .ZN(n286) );
  AOI31D0 U147 ( .A1(mantissa_ab[0]), .A2(n337), .A3(mantissa_c[0]), .B(n242), 
        .ZN(n295) );
  OAI21D0 U148 ( .A1(n338), .A2(n241), .B(n339), .ZN(n242) );
  AN2D0 U149 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .Z(n338) );
  CKND0 U150 ( .I(n241), .ZN(n337) );
  ND3D0 U151 ( .A1(mantissa_ab[2]), .A2(n339), .A3(mantissa_c[2]), .ZN(n241)
         );
  AN3D0 U152 ( .A1(n340), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .Z(n339) );
  OA211D0 U153 ( .A1(n341), .A2(n244), .B(n342), .C(n245), .Z(n218) );
  IAO21D0 U154 ( .A1(n246), .A2(n343), .B(n340), .ZN(n245) );
  AN3D0 U155 ( .A1(mantissa_ab[4]), .A2(n246), .A3(mantissa_c[4]), .Z(n340) );
  NR3D0 U156 ( .A1(n312), .A2(n343), .A3(n313), .ZN(n246) );
  CKND0 U157 ( .I(mantissa_c[5]), .ZN(n313) );
  IND4D0 U158 ( .A1(n244), .B1(mantissa_ab[6]), .B2(mantissa_ab[7]), .B3(n344), 
        .ZN(n343) );
  INR2D0 U159 ( .A1(mantissa_c[6]), .B1(n332), .ZN(n344) );
  CKND0 U160 ( .I(mantissa_ab[5]), .ZN(n312) );
  ND3D0 U161 ( .A1(mantissa_ab[8]), .A2(n342), .A3(mantissa_c[8]), .ZN(n244)
         );
  INR4D0 U162 ( .A1(n283), .B1(n334), .B2(n333), .B3(n206), .ZN(n342) );
  IND4D0 U163 ( .A1(n281), .B1(mantissa_ab[11]), .B2(mantissa_ab[12]), .B3(
        n345), .ZN(n206) );
  AN2D0 U164 ( .A1(mantissa_c[11]), .A2(mantissa_c[12]), .Z(n345) );
  ND3D0 U165 ( .A1(mantissa_ab[13]), .A2(n252), .A3(mantissa_c[13]), .ZN(n281)
         );
  NR2D0 U166 ( .A1(n280), .A2(n282), .ZN(n252) );
  CKND2D0 U167 ( .A1(mantissa_c[14]), .A2(mantissa_ab[14]), .ZN(n282) );
  ND4D0 U168 ( .A1(mantissa_ab[15]), .A2(n294), .A3(mantissa_ab[16]), .A4(n346), .ZN(n280) );
  NR2D0 U169 ( .A1(n335), .A2(n293), .ZN(n346) );
  CKND0 U170 ( .I(mantissa_c[16]), .ZN(n293) );
  CKND0 U171 ( .I(mantissa_c[15]), .ZN(n335) );
  CKND0 U172 ( .I(n204), .ZN(n294) );
  ND3D0 U173 ( .A1(mantissa_ab[17]), .A2(n290), .A3(mantissa_c[17]), .ZN(n204)
         );
  AN3D0 U174 ( .A1(n288), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .Z(n290)
         );
  NR4D0 U175 ( .A1(n261), .A2(n326), .A3(n325), .A4(n289), .ZN(n288) );
  CKND2D0 U176 ( .A1(mantissa_c[20]), .A2(mantissa_ab[20]), .ZN(n289) );
  CKND0 U177 ( .I(mantissa_ab[19]), .ZN(n325) );
  CKND0 U178 ( .I(mantissa_c[19]), .ZN(n326) );
  CKND2D0 U179 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .ZN(n261) );
  CKND0 U180 ( .I(mantissa_ab[9]), .ZN(n333) );
  CKND0 U181 ( .I(mantissa_c[9]), .ZN(n334) );
  AN2D0 U182 ( .A1(mantissa_c[10]), .A2(mantissa_ab[10]), .Z(n283) );
  NR2D0 U183 ( .A1(n331), .A2(n332), .ZN(n341) );
  CKND0 U184 ( .I(mantissa_c[7]), .ZN(n332) );
  CKND0 U185 ( .I(mantissa_ab[7]), .ZN(n331) );
  CKND0 U186 ( .I(sign_c), .ZN(n185) );
endmodule


module fma_aligner_adder_DW_rash_0_1 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108;

  MUX2ND0 U96 ( .I0(n106), .I1(n89), .S(n107), .ZN(n30) );
  AN3XD1 U54 ( .A1(SH[4]), .A2(n107), .A3(n108), .Z(n45) );
  OR2D1 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  OR2D1 U101 ( .A1(SH[4]), .A2(n108), .Z(n31) );
  NR2D1 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D1 U4 ( .A1(n103), .A2(SH[1]), .ZN(n52) );
  NR2D1 U5 ( .A1(n107), .A2(n31), .ZN(n36) );
  INVD1 U6 ( .I(n47), .ZN(n98) );
  NR2D1 U7 ( .A1(n27), .A2(n98), .ZN(B[17]) );
  NR2D1 U8 ( .A1(n50), .A2(n98), .ZN(B[19]) );
  NR2D1 U9 ( .A1(n58), .A2(n98), .ZN(B[18]) );
  OAI222D0 U10 ( .A1(n70), .A2(n26), .B1(n99), .B2(n61), .C1(n29), .C2(n98), 
        .ZN(B[12]) );
  NR2D1 U11 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D1 U12 ( .A1(n25), .A2(n98), .B1(n27), .B2(n26), .ZN(B[13]) );
  INVD1 U13 ( .I(n37), .ZN(n99) );
  NR2D1 U14 ( .A1(n98), .A2(n61), .ZN(B[20]) );
  INVD1 U15 ( .I(n58), .ZN(n87) );
  INVD1 U16 ( .I(n27), .ZN(n85) );
  INVD1 U17 ( .I(n59), .ZN(n91) );
  INVD1 U18 ( .I(n51), .ZN(n90) );
  INVD1 U19 ( .I(n25), .ZN(n92) );
  INVD1 U20 ( .I(n50), .ZN(n86) );
  INVD1 U21 ( .I(n70), .ZN(n89) );
  INVD1 U22 ( .I(n61), .ZN(n106) );
  AOI222D0 U23 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n102), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  IND2D1 U24 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  OAI211D1 U25 ( .A1(n29), .A2(n100), .B(n75), .C(n76), .ZN(B[0]) );
  INVD1 U26 ( .I(n36), .ZN(n100) );
  OA22D0 U27 ( .A1(n99), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  OAI222D0 U28 ( .A1(n59), .A2(n26), .B1(n58), .B2(n99), .C1(n38), .C2(n98), 
        .ZN(B[10]) );
  OAI22D1 U29 ( .A1(n59), .A2(n98), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI222D0 U30 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n98), 
        .ZN(B[8]) );
  OAI222D0 U31 ( .A1(n51), .A2(n26), .B1(n50), .B2(n99), .C1(n33), .C2(n98), 
        .ZN(B[11]) );
  OAI22D1 U32 ( .A1(n51), .A2(n98), .B1(n50), .B2(n26), .ZN(B[15]) );
  AOI221D0 U33 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U34 ( .A1(A[11]), .A2(n104), .B1(A[10]), .B2(n102), .Z(n78) );
  AOI221D0 U35 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29)
         );
  AO22D0 U36 ( .A1(A[15]), .A2(n104), .B1(A[14]), .B2(n102), .Z(n84) );
  AOI221D0 U37 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U38 ( .A1(A[12]), .A2(n104), .B1(A[11]), .B2(n102), .Z(n66) );
  AOI221D0 U39 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U40 ( .A1(A[20]), .A2(n104), .B1(A[19]), .B2(n102), .Z(n68) );
  AOI22D1 U41 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U42 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U43 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n102), .Z(n73) );
  AOI221D0 U44 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U45 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n102), .Z(n71) );
  AOI221D0 U46 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U47 ( .A1(A[17]), .A2(n104), .B1(A[16]), .B2(n102), .Z(n74) );
  AOI221D0 U48 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U49 ( .A1(A[18]), .A2(n104), .B1(A[17]), .B2(n102), .Z(n72) );
  AOI221D0 U50 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U51 ( .A1(A[16]), .A2(n104), .B1(A[15]), .B2(n102), .Z(n69) );
  AOI221D0 U52 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U53 ( .A1(A[19]), .A2(n104), .B1(A[18]), .B2(n102), .Z(n83) );
  OAI222D0 U55 ( .A1(n25), .A2(n26), .B1(n27), .B2(n99), .C1(n28), .C2(n98), 
        .ZN(B[9]) );
  NR2D1 U56 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  NR2D1 U57 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  ND2D1 U58 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  INVD1 U59 ( .I(n53), .ZN(n105) );
  INVD1 U60 ( .I(n52), .ZN(n101) );
  INVD1 U61 ( .I(n81), .ZN(n102) );
  INVD1 U62 ( .I(n80), .ZN(n104) );
  INVD1 U63 ( .I(SH[0]), .ZN(n103) );
  INVD1 U64 ( .I(SH[2]), .ZN(n107) );
  INVD1 U65 ( .I(SH[3]), .ZN(n108) );
  OAI221D0 U66 ( .A1(n28), .A2(n99), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U67 ( .A1(n36), .A2(n92), .B1(n45), .B2(n85), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U68 ( .A1(n101), .A2(n96), .B1(n105), .B2(n97), .C(n64), .ZN(n63)
         );
  OAI221D0 U69 ( .A1(n38), .A2(n99), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U70 ( .A1(n36), .A2(n91), .B1(n45), .B2(n87), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U71 ( .A1(n101), .A2(n95), .B1(n105), .B2(n96), .C(n57), .ZN(n56)
         );
  OAI221D0 U72 ( .A1(n33), .A2(n99), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U73 ( .A1(n36), .A2(n90), .B1(n45), .B2(n86), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U74 ( .A1(n101), .A2(n94), .B1(n105), .B2(n95), .C(n49), .ZN(n48)
         );
  OAI221D0 U75 ( .A1(n32), .A2(n26), .B1(n43), .B2(n98), .C(n44), .ZN(B[4]) );
  AOI222D0 U76 ( .A1(n37), .A2(n93), .B1(n45), .B2(n106), .C1(n36), .C2(n89), 
        .ZN(n44) );
  INVD1 U77 ( .I(n29), .ZN(n93) );
  OAI221D0 U78 ( .A1(n28), .A2(n26), .B1(n41), .B2(n98), .C(n42), .ZN(B[5]) );
  AOI22D1 U79 ( .A1(n36), .A2(n85), .B1(n37), .B2(n92), .ZN(n42) );
  OAI221D0 U80 ( .A1(n38), .A2(n26), .B1(n39), .B2(n98), .C(n40), .ZN(B[6]) );
  AOI22D1 U81 ( .A1(n36), .A2(n87), .B1(n37), .B2(n91), .ZN(n40) );
  OAI221D0 U82 ( .A1(n33), .A2(n26), .B1(n34), .B2(n98), .C(n35), .ZN(B[7]) );
  AOI22D1 U83 ( .A1(n36), .A2(n86), .B1(n37), .B2(n90), .ZN(n35) );
  AOI221D0 U84 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U85 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n102), .Z(n54) );
  AOI221D0 U86 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U87 ( .A1(A[7]), .A2(n104), .B1(A[6]), .B2(n102), .Z(n77) );
  AOI221D0 U88 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U89 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n102), .Z(n60) );
  AOI221D0 U90 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U91 ( .A1(A[8]), .A2(n104), .B1(A[7]), .B2(n102), .Z(n65) );
  AOI22D1 U92 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n102), .ZN(n57) );
  AOI22D1 U93 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n102), .ZN(n49) );
  AOI22D1 U94 ( .A1(A[4]), .A2(n104), .B1(A[3]), .B2(n102), .ZN(n64) );
  ND2D1 U97 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  ND2D1 U98 ( .A1(SH[1]), .A2(n103), .ZN(n81) );
  AOI32D1 U99 ( .A1(n88), .A2(n108), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75)
         );
  INVD1 U100 ( .I(n30), .ZN(n88) );
  OAI221D0 U102 ( .A1(n80), .A2(n95), .B1(n81), .B2(n96), .C(n82), .ZN(n79) );
  AOI22D1 U103 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  INVD1 U104 ( .I(A[4]), .ZN(n94) );
  INVD1 U105 ( .I(A[3]), .ZN(n95) );
  INVD1 U106 ( .I(A[2]), .ZN(n96) );
  INVD1 U107 ( .I(A[1]), .ZN(n97) );
endmodule


module fma_aligner_adder_1 ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n633, n634, n658,
         n848, n850, n872, n905, n906, n946, n951, n1063, n1103, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;
  assign mantissa_ab_c[21] = n1147;

  CKXOR2D1 U1204 ( .A1(n850), .A2(n872), .Z(n545) );
  CKXOR2D1 U1205 ( .A1(n532), .A2(n545), .Z(n848) );
  CKXOR2D1 U1206 ( .A1(n633), .A2(n634), .Z(n536) );
  CKXOR2D1 U1207 ( .A1(n946), .A2(n531), .Z(n546) );
  CKXOR2D1 U1208 ( .A1(n1103), .A2(n543), .Z(n547) );
  CKXOR2D1 U1209 ( .A1(n546), .A2(n547), .Z(n634) );
  CKXOR2D1 U1210 ( .A1(n658), .A2(n537), .Z(n538) );
  CKXOR2D1 U1211 ( .A1(n951), .A2(n529), .Z(n548) );
  CKXOR2D1 U1212 ( .A1(n542), .A2(n530), .Z(n549) );
  CKXOR2D1 U1213 ( .A1(n548), .A2(n549), .Z(n537) );
  CKXOR2D1 U1214 ( .A1(n540), .A2(n539), .Z(n541) );
  CKXOR2D1 U1215 ( .A1(n905), .A2(n906), .Z(n550) );
  CKXOR2D1 U1216 ( .A1(n1063), .A2(n544), .Z(n551) );
  CKXOR2D1 U1217 ( .A1(n550), .A2(n551), .Z(n539) );
  fma_lza_1 fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0_1 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(
        n552), .SH(exp_diff), .SH_TC(n552), .B({N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45}) );
  TIEL U600 ( .ZN(n552) );
  OAI21D0 U601 ( .A1(n1), .A2(n2), .B(n3), .ZN(sign_ab_c) );
  MUX2ND0 U602 ( .I0(n4), .I1(c[15]), .S(fma_byp), .ZN(n3) );
  AOI31D0 U603 ( .A1(n5), .A2(n6), .A3(n7), .B(n8), .ZN(n4) );
  OAI21D0 U604 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  CKND0 U605 ( .I(exp_ab_less), .ZN(n11) );
  OA31D0 U606 ( .A1(n10), .A2(exp_ab_greater), .A3(n9), .B(n12), .Z(n1) );
  NR2D0 U607 ( .A1(n13), .A2(c[9]), .ZN(n9) );
  OA221D0 U608 ( .A1(mantissa_ab[8]), .A2(n14), .B1(mantissa_ab[9]), .B2(n15), 
        .C(n16), .Z(n10) );
  AO22D0 U609 ( .A1(n14), .A2(mantissa_ab[8]), .B1(n17), .B2(n18), .Z(n16) );
  OAI221D0 U610 ( .A1(c[7]), .A2(n19), .B1(c[6]), .B2(n20), .C(n21), .ZN(n18)
         );
  OAI222D0 U611 ( .A1(mantissa_ab[5]), .A2(n22), .B1(mantissa_ab[6]), .B2(n23), 
        .C1(n24), .C2(n25), .ZN(n21) );
  MAOI222D0 U612 ( .A(n26), .B(n27), .C(c[4]), .ZN(n25) );
  AOI22D0 U613 ( .A1(mantissa_ab[3]), .A2(n28), .B1(n29), .B2(n30), .ZN(n27)
         );
  OR2D0 U614 ( .A1(n29), .A2(n30), .Z(n28) );
  MAOI22D0 U615 ( .A1(n31), .A2(c[2]), .B1(mantissa_ab[2]), .B2(n32), .ZN(n29)
         );
  NR2D0 U616 ( .A1(c[2]), .A2(n31), .ZN(n32) );
  OAI22D0 U617 ( .A1(n33), .A2(n34), .B1(mantissa_ab[1]), .B2(n35), .ZN(n31)
         );
  INR2D0 U618 ( .A1(n33), .B1(c[1]), .ZN(n35) );
  NR2D0 U619 ( .A1(n36), .A2(c[0]), .ZN(n33) );
  NR2D0 U620 ( .A1(c[5]), .A2(n37), .ZN(n24) );
  CKND2D0 U621 ( .A1(c[7]), .A2(n19), .ZN(n17) );
  AOI31D0 U622 ( .A1(n38), .A2(n39), .A3(n40), .B(n41), .ZN(n658) );
  OAI21D0 U623 ( .A1(n42), .A2(n43), .B(n44), .ZN(n39) );
  AOI21D0 U624 ( .A1(n45), .A2(n46), .B(n47), .ZN(n42) );
  AOI21D0 U625 ( .A1(n537), .A2(n48), .B(n49), .ZN(n633) );
  IOA21D0 U626 ( .A1(n50), .A2(n38), .B(n51), .ZN(n48) );
  CKND0 U627 ( .I(n52), .ZN(n540) );
  NR3D0 U628 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1147) );
  MUX2ND0 U629 ( .I0(n56), .I1(n57), .S(n58), .ZN(mantissa_ab_c[9]) );
  IAO21D0 U630 ( .A1(n59), .A2(fma_byp), .B(n60), .ZN(n57) );
  CKND2D0 U631 ( .A1(n61), .A2(n59), .ZN(n56) );
  MUX2ND0 U632 ( .I0(n62), .I1(n63), .S(n64), .ZN(mantissa_ab_c[8]) );
  CKND2D0 U633 ( .A1(n61), .A2(n65), .ZN(n63) );
  IAO21D0 U634 ( .A1(n65), .A2(fma_byp), .B(n60), .ZN(n62) );
  MUX2ND0 U635 ( .I0(n66), .I1(n67), .S(n68), .ZN(mantissa_ab_c[7]) );
  CKND2D0 U636 ( .A1(n61), .A2(n69), .ZN(n67) );
  AOI21D0 U637 ( .A1(n70), .A2(n71), .B(n60), .ZN(n66) );
  MUX2ND0 U638 ( .I0(n72), .I1(n73), .S(n74), .ZN(mantissa_ab_c[6]) );
  OR2D0 U639 ( .A1(n75), .A2(n53), .Z(n73) );
  AOI21D0 U640 ( .A1(n75), .A2(n71), .B(n60), .ZN(n72) );
  MUX2ND0 U641 ( .I0(n76), .I1(n77), .S(n78), .ZN(mantissa_ab_c[5]) );
  CKND2D0 U642 ( .A1(n61), .A2(n79), .ZN(n77) );
  IAO21D0 U643 ( .A1(n79), .A2(fma_byp), .B(n60), .ZN(n76) );
  MUX2ND0 U644 ( .I0(n80), .I1(n81), .S(n82), .ZN(mantissa_ab_c[4]) );
  IND2D0 U645 ( .A1(n83), .B1(n61), .ZN(n81) );
  AOI21D0 U646 ( .A1(n83), .A2(n71), .B(n60), .ZN(n80) );
  MUX2ND0 U647 ( .I0(n84), .I1(n85), .S(n86), .ZN(mantissa_ab_c[3]) );
  CKND2D0 U648 ( .A1(n61), .A2(n87), .ZN(n85) );
  IAO21D0 U649 ( .A1(n87), .A2(fma_byp), .B(n60), .ZN(n84) );
  MUX2ND0 U650 ( .I0(n88), .I1(n89), .S(n90), .ZN(mantissa_ab_c[2]) );
  OR2D0 U651 ( .A1(n91), .A2(n53), .Z(n89) );
  AOI21D0 U652 ( .A1(n91), .A2(n71), .B(n60), .ZN(n88) );
  OAI21D0 U653 ( .A1(n92), .A2(n71), .B(n93), .ZN(mantissa_ab_c[20]) );
  MUX2ND0 U654 ( .I0(n94), .I1(n95), .S(n55), .ZN(n93) );
  MUX2ND0 U655 ( .I0(n96), .I1(n536), .S(n5), .ZN(n55) );
  OAI21D0 U656 ( .A1(fma_byp), .A2(n54), .B(n97), .ZN(n95) );
  INR2D0 U657 ( .A1(n54), .B1(n53), .ZN(n94) );
  CKND2D0 U658 ( .A1(n98), .A2(n99), .ZN(n54) );
  MUX2ND0 U659 ( .I0(n100), .I1(n101), .S(n102), .ZN(mantissa_ab_c[1]) );
  AOI21D0 U660 ( .A1(n103), .A2(n71), .B(n60), .ZN(n101) );
  CKND2D0 U661 ( .A1(n104), .A2(n61), .ZN(n100) );
  CKND0 U662 ( .I(n53), .ZN(n61) );
  OAI21D0 U663 ( .A1(n15), .A2(n71), .B(n105), .ZN(mantissa_ab_c[19]) );
  MUX2ND0 U664 ( .I0(n106), .I1(n107), .S(n99), .ZN(n105) );
  MUX2D0 U665 ( .I0(n108), .I1(n538), .S(n5), .Z(n99) );
  NR2D0 U666 ( .A1(n98), .A2(n53), .ZN(n107) );
  CKND0 U667 ( .I(n109), .ZN(n98) );
  OAI21D0 U668 ( .A1(fma_byp), .A2(n109), .B(n97), .ZN(n106) );
  CKND2D0 U669 ( .A1(n110), .A2(n111), .ZN(n109) );
  OAI21D0 U670 ( .A1(n14), .A2(n71), .B(n112), .ZN(mantissa_ab_c[18]) );
  MUX2ND0 U671 ( .I0(n113), .I1(n114), .S(n111), .ZN(n112) );
  MUX2ND0 U672 ( .I0(n115), .I1(n116), .S(add_byp), .ZN(n111) );
  CKXOR2D0 U673 ( .A1(n38), .A2(n50), .Z(n115) );
  OAI221D0 U674 ( .A1(n117), .A2(n44), .B1(n117), .B2(n118), .C(n119), .ZN(n50) );
  IND2D0 U675 ( .A1(n43), .B1(n120), .ZN(n118) );
  NR2D0 U676 ( .A1(n110), .A2(n53), .ZN(n114) );
  CKND0 U677 ( .I(n121), .ZN(n110) );
  OAI21D0 U678 ( .A1(fma_byp), .A2(n121), .B(n97), .ZN(n113) );
  CKND2D0 U679 ( .A1(n122), .A2(n123), .ZN(n121) );
  OAI21D0 U680 ( .A1(n124), .A2(n71), .B(n125), .ZN(mantissa_ab_c[17]) );
  MUX2ND0 U681 ( .I0(n126), .I1(n127), .S(n123), .ZN(n125) );
  MUX2ND0 U682 ( .I0(n128), .I1(n129), .S(add_byp), .ZN(n123) );
  CKXOR2D0 U683 ( .A1(n130), .A2(n40), .Z(n128) );
  NR2D0 U684 ( .A1(n122), .A2(n53), .ZN(n127) );
  CKND0 U685 ( .I(n131), .ZN(n122) );
  OAI21D0 U686 ( .A1(fma_byp), .A2(n131), .B(n97), .ZN(n126) );
  CKND2D0 U687 ( .A1(n132), .A2(n133), .ZN(n131) );
  OAI21D0 U688 ( .A1(n23), .A2(n71), .B(n134), .ZN(mantissa_ab_c[16]) );
  MUX2ND0 U689 ( .I0(n135), .I1(n136), .S(n133), .ZN(n134) );
  MUX2ND0 U690 ( .I0(n137), .I1(n138), .S(add_byp), .ZN(n133) );
  XNR2D0 U691 ( .A1(n120), .A2(n43), .ZN(n137) );
  OAI21D0 U692 ( .A1(n139), .A2(n140), .B(n141), .ZN(n120) );
  NR2D0 U693 ( .A1(n132), .A2(n53), .ZN(n136) );
  CKND0 U694 ( .I(n142), .ZN(n132) );
  OAI21D0 U695 ( .A1(fma_byp), .A2(n142), .B(n97), .ZN(n135) );
  CKND2D0 U696 ( .A1(n143), .A2(n144), .ZN(n142) );
  OAI21D0 U697 ( .A1(n22), .A2(n71), .B(n145), .ZN(mantissa_ab_c[15]) );
  MUX2ND0 U698 ( .I0(n146), .I1(n147), .S(n144), .ZN(n145) );
  MUX2D0 U699 ( .I0(n148), .I1(n149), .S(n5), .Z(n144) );
  CKXOR2D0 U700 ( .A1(n46), .A2(n139), .Z(n149) );
  CKND2D0 U701 ( .A1(n150), .A2(n140), .ZN(n46) );
  NR2D0 U702 ( .A1(n143), .A2(n53), .ZN(n147) );
  CKND0 U703 ( .I(n151), .ZN(n143) );
  OAI21D0 U704 ( .A1(fma_byp), .A2(n151), .B(n97), .ZN(n146) );
  CKND2D0 U705 ( .A1(n152), .A2(n153), .ZN(n151) );
  OAI21D0 U706 ( .A1(n154), .A2(n71), .B(n155), .ZN(mantissa_ab_c[14]) );
  MUX2ND0 U707 ( .I0(n156), .I1(n157), .S(n153), .ZN(n155) );
  MUX2D0 U708 ( .I0(n158), .I1(n159), .S(n5), .Z(n153) );
  OAI21D0 U709 ( .A1(n160), .A2(n161), .B(n140), .ZN(n159) );
  CKND2D0 U710 ( .A1(n160), .A2(n161), .ZN(n140) );
  OAI221D0 U711 ( .A1(n162), .A2(n163), .B1(n162), .B2(n164), .C(n165), .ZN(
        n161) );
  NR2D0 U712 ( .A1(n152), .A2(n53), .ZN(n157) );
  CKND0 U713 ( .I(n166), .ZN(n152) );
  OAI21D0 U714 ( .A1(fma_byp), .A2(n166), .B(n97), .ZN(n156) );
  CKND2D0 U715 ( .A1(n167), .A2(n168), .ZN(n166) );
  OAI21D0 U716 ( .A1(n30), .A2(n71), .B(n169), .ZN(mantissa_ab_c[13]) );
  MUX2ND0 U717 ( .I0(n170), .I1(n171), .S(n168), .ZN(n169) );
  MUX2ND0 U718 ( .I0(n172), .I1(n173), .S(add_byp), .ZN(n168) );
  CKXOR2D0 U719 ( .A1(n162), .A2(n174), .Z(n172) );
  NR2D0 U720 ( .A1(n167), .A2(n53), .ZN(n171) );
  CKND0 U721 ( .I(n175), .ZN(n167) );
  OAI21D0 U722 ( .A1(fma_byp), .A2(n175), .B(n97), .ZN(n170) );
  CKND2D0 U723 ( .A1(n176), .A2(n177), .ZN(n175) );
  OAI21D0 U724 ( .A1(n178), .A2(n71), .B(n179), .ZN(mantissa_ab_c[12]) );
  MUX2ND0 U725 ( .I0(n180), .I1(n181), .S(n177), .ZN(n179) );
  MUX2ND0 U726 ( .I0(n182), .I1(n183), .S(add_byp), .ZN(n177) );
  OA21D0 U727 ( .A1(n184), .A2(n185), .B(n164), .Z(n182) );
  NR2D0 U728 ( .A1(n176), .A2(n53), .ZN(n181) );
  CKND0 U729 ( .I(n186), .ZN(n176) );
  OAI21D0 U730 ( .A1(fma_byp), .A2(n186), .B(n97), .ZN(n180) );
  CKND2D0 U731 ( .A1(n187), .A2(n188), .ZN(n186) );
  OAI21D0 U732 ( .A1(n34), .A2(n71), .B(n189), .ZN(mantissa_ab_c[11]) );
  MUX2ND0 U733 ( .I0(n190), .I1(n191), .S(n188), .ZN(n189) );
  MUX2D0 U734 ( .I0(n192), .I1(n193), .S(n5), .Z(n188) );
  OAI21D0 U735 ( .A1(n194), .A2(n195), .B(n196), .ZN(n193) );
  NR2D0 U736 ( .A1(n187), .A2(n53), .ZN(n191) );
  CKND0 U737 ( .I(n197), .ZN(n187) );
  OAI21D0 U738 ( .A1(fma_byp), .A2(n197), .B(n97), .ZN(n190) );
  CKND2D0 U739 ( .A1(n198), .A2(n199), .ZN(n197) );
  OAI21D0 U740 ( .A1(n71), .A2(n200), .B(n201), .ZN(mantissa_ab_c[10]) );
  MUX2ND0 U741 ( .I0(n202), .I1(n203), .S(n199), .ZN(n201) );
  MUX2ND0 U742 ( .I0(n204), .I1(n205), .S(add_byp), .ZN(n199) );
  CKXOR2D0 U743 ( .A1(n206), .A2(n207), .Z(n204) );
  NR2D0 U744 ( .A1(n198), .A2(n53), .ZN(n203) );
  CKND2D0 U745 ( .A1(n208), .A2(n71), .ZN(n53) );
  CKXOR2D0 U746 ( .A1(n209), .A2(n210), .Z(n208) );
  AO21D0 U747 ( .A1(n71), .A2(n198), .B(n60), .Z(n202) );
  CKND0 U748 ( .I(n97), .ZN(n60) );
  MUX2ND0 U749 ( .I0(comp_mantissa_ab[21]), .I1(n211), .S(n210), .ZN(n97) );
  CKND2D0 U750 ( .A1(n212), .A2(n5), .ZN(n210) );
  CKXOR2D0 U751 ( .A1(n213), .A2(n214), .Z(n212) );
  MAOI22D0 U752 ( .A1(n634), .A2(n215), .B1(n216), .B2(n96), .ZN(n213) );
  AO21D0 U753 ( .A1(n217), .A2(n537), .B(n49), .Z(n215) );
  NR2D0 U754 ( .A1(n108), .A2(n218), .ZN(n49) );
  AO31D0 U755 ( .A1(n38), .A2(n130), .A3(n40), .B(n41), .Z(n217) );
  OAI21D0 U756 ( .A1(n219), .A2(n119), .B(n51), .ZN(n41) );
  CKND0 U757 ( .I(n117), .ZN(n40) );
  OAI21D0 U758 ( .A1(n129), .A2(n220), .B(n119), .ZN(n117) );
  CKND2D0 U759 ( .A1(n129), .A2(n220), .ZN(n119) );
  OAI21D0 U760 ( .A1(n221), .A2(n43), .B(n44), .ZN(n130) );
  OAI21D0 U761 ( .A1(n138), .A2(n222), .B(n44), .ZN(n43) );
  CKND2D0 U762 ( .A1(n138), .A2(n222), .ZN(n44) );
  AOI31D0 U763 ( .A1(n160), .A2(n223), .A3(n45), .B(n224), .ZN(n221) );
  CKND0 U764 ( .I(n141), .ZN(n224) );
  IAO21D0 U765 ( .A1(n139), .A2(n150), .B(n47), .ZN(n141) );
  CKND0 U766 ( .I(n45), .ZN(n139) );
  AOI21D0 U767 ( .A1(n225), .A2(n148), .B(n47), .ZN(n45) );
  NR2D0 U768 ( .A1(n148), .A2(n225), .ZN(n47) );
  OAI21D0 U769 ( .A1(n174), .A2(n162), .B(n165), .ZN(n223) );
  OAI21D0 U770 ( .A1(n226), .A2(n173), .B(n165), .ZN(n162) );
  CKND2D0 U771 ( .A1(n226), .A2(n173), .ZN(n165) );
  CKND0 U772 ( .I(n227), .ZN(n226) );
  AN2D0 U773 ( .A1(n164), .A2(n163), .Z(n174) );
  CKND2D0 U774 ( .A1(n184), .A2(n185), .ZN(n164) );
  OAI21D0 U775 ( .A1(n192), .A2(n228), .B(n196), .ZN(n185) );
  CKND2D0 U776 ( .A1(n194), .A2(n195), .ZN(n196) );
  OAI21D0 U777 ( .A1(n206), .A2(n207), .B(n229), .ZN(n195) );
  OAI21D0 U778 ( .A1(n230), .A2(n205), .B(n229), .ZN(n207) );
  CKND2D0 U779 ( .A1(n205), .A2(n230), .ZN(n229) );
  MAOI22D0 U780 ( .A1(n539), .A2(n52), .B1(n231), .B2(n232), .ZN(n206) );
  OAI21D0 U781 ( .A1(n233), .A2(n234), .B(n235), .ZN(n52) );
  CKXOR2D0 U782 ( .A1(n192), .A2(n228), .Z(n194) );
  OA21D0 U783 ( .A1(n236), .A2(n183), .B(n163), .Z(n184) );
  CKND2D0 U784 ( .A1(n236), .A2(n183), .ZN(n163) );
  CKND0 U785 ( .I(n237), .ZN(n236) );
  OA21D0 U786 ( .A1(n238), .A2(n239), .B(n150), .Z(n160) );
  CKND2D0 U787 ( .A1(n238), .A2(n239), .ZN(n150) );
  CKND0 U788 ( .I(n240), .ZN(n239) );
  CKND0 U789 ( .I(n219), .ZN(n38) );
  OAI21D0 U790 ( .A1(n116), .A2(n241), .B(n51), .ZN(n219) );
  CKND2D0 U791 ( .A1(n116), .A2(n241), .ZN(n51) );
  CKND0 U792 ( .I(n242), .ZN(n241) );
  AN2D0 U793 ( .A1(n209), .A2(n71), .Z(n211) );
  NR2D0 U794 ( .A1(n59), .A2(n58), .ZN(n198) );
  MUX2ND0 U795 ( .I0(n541), .I1(n231), .S(add_byp), .ZN(n58) );
  IND2D0 U796 ( .A1(n65), .B1(n64), .ZN(n59) );
  MUX2ND0 U797 ( .I0(n243), .I1(n244), .S(add_byp), .ZN(n64) );
  CKXOR2D0 U798 ( .A1(n234), .A2(n233), .Z(n243) );
  OA22D0 U799 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .Z(n233) );
  OAI21D0 U800 ( .A1(n249), .A2(n244), .B(n235), .ZN(n234) );
  CKND2D0 U801 ( .A1(n244), .A2(n249), .ZN(n235) );
  CKND0 U802 ( .I(n250), .ZN(n249) );
  CKND2D0 U803 ( .A1(n70), .A2(n68), .ZN(n65) );
  MUX2D0 U804 ( .I0(n245), .I1(n251), .S(n5), .Z(n68) );
  XNR2D0 U805 ( .A1(n247), .A2(n248), .ZN(n251) );
  XNR2D0 U806 ( .A1(n245), .A2(n246), .ZN(n248) );
  OA21D0 U807 ( .A1(n252), .A2(n253), .B(n254), .Z(n247) );
  CKND0 U808 ( .I(n69), .ZN(n70) );
  CKND2D0 U809 ( .A1(n75), .A2(n74), .ZN(n69) );
  MUX2D0 U810 ( .I0(n255), .I1(n256), .S(n5), .Z(n74) );
  XNR2D0 U811 ( .A1(n253), .A2(n252), .ZN(n256) );
  AOI21D0 U812 ( .A1(n257), .A2(n258), .B(n259), .ZN(n252) );
  OAI21D0 U813 ( .A1(n260), .A2(n261), .B(n254), .ZN(n253) );
  CKND2D0 U814 ( .A1(n260), .A2(n261), .ZN(n254) );
  CKND0 U815 ( .I(n255), .ZN(n260) );
  INR2D0 U816 ( .A1(n78), .B1(n79), .ZN(n75) );
  CKND2D0 U817 ( .A1(n83), .A2(n82), .ZN(n79) );
  MUX2ND0 U818 ( .I0(n262), .I1(n263), .S(add_byp), .ZN(n82) );
  CKXOR2D0 U819 ( .A1(n264), .A2(n265), .Z(n262) );
  INR2D0 U820 ( .A1(n86), .B1(n87), .ZN(n83) );
  CKND2D0 U821 ( .A1(n91), .A2(n90), .ZN(n87) );
  MUX2ND0 U822 ( .I0(n266), .I1(n267), .S(add_byp), .ZN(n90) );
  OA21D0 U823 ( .A1(n268), .A2(n269), .B(n270), .Z(n266) );
  NR2D0 U824 ( .A1(n102), .A2(n104), .ZN(n91) );
  CKXOR2D0 U825 ( .A1(n271), .A2(n272), .Z(n102) );
  CKND2D0 U826 ( .A1(n848), .A2(n5), .ZN(n272) );
  MUX2ND0 U827 ( .I0(n273), .I1(n274), .S(add_byp), .ZN(n86) );
  CKXOR2D0 U828 ( .A1(n275), .A2(n276), .Z(n273) );
  OAI22D0 U829 ( .A1(add_byp), .A2(n277), .B1(n257), .B2(n278), .ZN(n78) );
  AOI21D0 U830 ( .A1(n279), .A2(n280), .B(add_byp), .ZN(n278) );
  AOI31D0 U831 ( .A1(n258), .A2(n257), .A3(n279), .B(n259), .ZN(n277) );
  INR2D0 U832 ( .A1(n281), .B1(n279), .ZN(n259) );
  CKXOR2D0 U833 ( .A1(n280), .A2(n282), .Z(n281) );
  OA21D0 U834 ( .A1(n264), .A2(n265), .B(n283), .Z(n279) );
  OAI21D0 U835 ( .A1(n263), .A2(n284), .B(n283), .ZN(n265) );
  CKND2D0 U836 ( .A1(n263), .A2(n284), .ZN(n283) );
  CKND0 U837 ( .I(n285), .ZN(n263) );
  OA21D0 U838 ( .A1(n275), .A2(n276), .B(n286), .Z(n264) );
  OAI21D0 U839 ( .A1(n274), .A2(n287), .B(n286), .ZN(n276) );
  CKND2D0 U840 ( .A1(n274), .A2(n287), .ZN(n286) );
  CKND0 U841 ( .I(n288), .ZN(n287) );
  AN2D0 U842 ( .A1(n270), .A2(n289), .Z(n275) );
  CKND2D0 U843 ( .A1(n268), .A2(n269), .ZN(n270) );
  OA21D0 U844 ( .A1(n267), .A2(n290), .B(n289), .Z(n269) );
  CKND2D0 U845 ( .A1(n267), .A2(n290), .ZN(n289) );
  CKND0 U846 ( .I(n291), .ZN(n268) );
  MAOI222D0 U847 ( .A(n292), .B(n850), .C(n293), .ZN(n291) );
  MUX2ND0 U848 ( .I0(n294), .I1(n295), .S(n296), .ZN(n293) );
  NR2D0 U849 ( .A1(n8), .A2(n297), .ZN(n294) );
  NR2D0 U850 ( .A1(n298), .A2(n297), .ZN(n850) );
  CKXOR2D0 U851 ( .A1(n872), .A2(n532), .Z(n292) );
  CKND0 U852 ( .I(n282), .ZN(n257) );
  CKND0 U853 ( .I(n280), .ZN(n258) );
  NR2D0 U854 ( .A1(fma_byp), .A2(n103), .ZN(mantissa_ab_c[0]) );
  CKND0 U855 ( .I(n104), .ZN(n103) );
  XNR2D0 U856 ( .A1(n299), .A2(n297), .ZN(n104) );
  MUX2D0 U857 ( .I0(c[14]), .I1(exp_ab[4]), .S(n300), .Z(exp_ab_c[4]) );
  MUX2D0 U858 ( .I0(c[13]), .I1(exp_ab[3]), .S(n300), .Z(exp_ab_c[3]) );
  MUX2ND0 U859 ( .I0(n301), .I1(n302), .S(n300), .ZN(exp_ab_c[2]) );
  MUX2ND0 U860 ( .I0(n303), .I1(n304), .S(n300), .ZN(exp_ab_c[1]) );
  MUX2ND0 U861 ( .I0(n305), .I1(n306), .S(n300), .ZN(exp_ab_c[0]) );
  NR2D0 U862 ( .A1(fma_byp), .A2(n307), .ZN(n300) );
  NR2D0 U863 ( .A1(fma_byp), .A2(n232), .ZN(comp_mantissa_c[9]) );
  CKXOR2D0 U864 ( .A1(n905), .A2(n308), .Z(n232) );
  CKND0 U865 ( .I(n309), .ZN(n905) );
  NR2D0 U866 ( .A1(fma_byp), .A2(n250), .ZN(comp_mantissa_c[8]) );
  CKND2D0 U867 ( .A1(n310), .A2(n311), .ZN(n250) );
  MUX2ND0 U868 ( .I0(n312), .I1(n313), .S(n314), .ZN(n310) );
  NR2D0 U869 ( .A1(n315), .A2(n312), .ZN(n313) );
  NR2D0 U870 ( .A1(fma_byp), .A2(n246), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U871 ( .A1(n316), .A2(n317), .ZN(n246) );
  MUX2ND0 U872 ( .I0(n318), .I1(n319), .S(n314), .ZN(n316) );
  NR2D0 U873 ( .A1(n320), .A2(n318), .ZN(n319) );
  INR2D0 U874 ( .A1(n261), .B1(fma_byp), .ZN(comp_mantissa_c[6]) );
  INR2D0 U875 ( .A1(n321), .B1(n320), .ZN(n261) );
  MUX2ND0 U876 ( .I0(n322), .I1(n323), .S(n314), .ZN(n321) );
  INR2D0 U877 ( .A1(n324), .B1(n322), .ZN(n323) );
  CKND0 U878 ( .I(n325), .ZN(n322) );
  NR2D0 U879 ( .A1(fma_byp), .A2(n280), .ZN(comp_mantissa_c[5]) );
  CKND2D0 U880 ( .A1(n326), .A2(n324), .ZN(n280) );
  MUX2ND0 U881 ( .I0(n327), .I1(n328), .S(n314), .ZN(n326) );
  NR2D0 U882 ( .A1(n327), .A2(n329), .ZN(n328) );
  CKND0 U883 ( .I(n330), .ZN(n327) );
  INR2D0 U884 ( .A1(n284), .B1(fma_byp), .ZN(comp_mantissa_c[4]) );
  INR3D0 U885 ( .A1(n331), .B1(n6), .B2(n329), .ZN(n284) );
  NR2D0 U886 ( .A1(n332), .A2(n333), .ZN(n329) );
  MUX2ND0 U887 ( .I0(n334), .I1(n335), .S(n314), .ZN(n331) );
  NR2D0 U888 ( .A1(n336), .A2(n334), .ZN(n335) );
  CKND0 U889 ( .I(n333), .ZN(n334) );
  NR2D0 U890 ( .A1(fma_byp), .A2(n288), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U891 ( .A1(n337), .A2(n332), .ZN(n288) );
  MUX2ND0 U892 ( .I0(n338), .I1(n339), .S(n314), .ZN(n337) );
  NR2D0 U893 ( .A1(n338), .A2(n340), .ZN(n339) );
  INR2D0 U894 ( .A1(n290), .B1(fma_byp), .ZN(comp_mantissa_c[2]) );
  INR2D0 U895 ( .A1(n341), .B1(n340), .ZN(n290) );
  MUX2ND0 U896 ( .I0(n2), .I1(n342), .S(n343), .ZN(n341) );
  OAI21D0 U897 ( .A1(n2), .A2(n344), .B(n345), .ZN(n342) );
  NR2D0 U898 ( .A1(fma_byp), .A2(n214), .ZN(comp_mantissa_c[21]) );
  CKND2D0 U899 ( .A1(n314), .A2(n346), .ZN(n214) );
  IND4D0 U900 ( .A1(n543), .B1(n347), .B2(n348), .B3(n349), .ZN(n346) );
  MUX2ND0 U901 ( .I0(n216), .I1(n92), .S(fma_byp), .ZN(comp_mantissa_c[20]) );
  XNR2D0 U902 ( .A1(n946), .A2(n543), .ZN(n216) );
  AOI211D0 U903 ( .A1(n350), .A2(exp_ab_greater), .B(n351), .C(n92), .ZN(n543)
         );
  AO21D0 U904 ( .A1(n314), .A2(n542), .B(n951), .Z(n946) );
  NR2D0 U905 ( .A1(fma_byp), .A2(n352), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U906 ( .A1(n872), .A2(n344), .Z(n352) );
  CKND0 U907 ( .I(n345), .ZN(n872) );
  CKND2D0 U908 ( .A1(n299), .A2(c[15]), .ZN(n345) );
  NR2D0 U909 ( .A1(n298), .A2(add_byp), .ZN(n299) );
  MUX2ND0 U910 ( .I0(n218), .I1(n15), .S(fma_byp), .ZN(comp_mantissa_c[19]) );
  XNR2D0 U911 ( .A1(n951), .A2(n542), .ZN(n218) );
  CKND0 U912 ( .I(n349), .ZN(n542) );
  CKND2D0 U913 ( .A1(n353), .A2(n354), .ZN(n349) );
  MUX2ND0 U914 ( .I0(n15), .I1(n355), .S(exp_ab_greater), .ZN(n353) );
  AOI21D0 U915 ( .A1(n348), .A2(n347), .B(n2), .ZN(n951) );
  MUX2ND0 U916 ( .I0(n242), .I1(n14), .S(fma_byp), .ZN(comp_mantissa_c[18]) );
  MUX2ND0 U917 ( .I0(n356), .I1(n357), .S(n348), .ZN(n242) );
  CKND2D0 U918 ( .A1(n358), .A2(n354), .ZN(n348) );
  MUX2ND0 U919 ( .I0(n14), .I1(n359), .S(exp_ab_greater), .ZN(n358) );
  OAI21D0 U920 ( .A1(n2), .A2(n360), .B(n361), .ZN(n357) );
  OR2D0 U921 ( .A1(n347), .A2(n2), .Z(n356) );
  INR3D0 U922 ( .A1(n360), .B1(n362), .B2(n363), .ZN(n347) );
  MUX2D0 U923 ( .I0(c[7]), .I1(n220), .S(n71), .Z(comp_mantissa_c[17]) );
  CKXOR2D0 U924 ( .A1(n361), .A2(n360), .Z(n220) );
  CKND2D0 U925 ( .A1(n364), .A2(n354), .ZN(n360) );
  MUX2ND0 U926 ( .I0(n124), .I1(n365), .S(exp_ab_greater), .ZN(n364) );
  OAI21D0 U927 ( .A1(n362), .A2(n363), .B(n314), .ZN(n361) );
  MUX2D0 U928 ( .I0(c[6]), .I1(n222), .S(n71), .Z(comp_mantissa_c[16]) );
  XNR2D0 U929 ( .A1(n362), .A2(n366), .ZN(n222) );
  CKND2D0 U930 ( .A1(n314), .A2(n363), .ZN(n366) );
  MUX2D0 U931 ( .I0(n367), .I1(c[6]), .S(n6), .Z(n362) );
  NR3D0 U932 ( .A1(n368), .A2(exp_diff[4]), .A3(exp_diff[3]), .ZN(n367) );
  MUX2ND0 U933 ( .I0(n225), .I1(n22), .S(fma_byp), .ZN(comp_mantissa_c[15]) );
  CKND2D0 U934 ( .A1(n369), .A2(n363), .ZN(n225) );
  CKND2D0 U935 ( .A1(n370), .A2(n371), .ZN(n363) );
  MUX2ND0 U936 ( .I0(n371), .I1(n372), .S(n314), .ZN(n369) );
  NR2D0 U937 ( .A1(n370), .A2(n371), .ZN(n372) );
  CKND0 U938 ( .I(n373), .ZN(n370) );
  MUX2D0 U939 ( .I0(n374), .I1(n22), .S(n6), .Z(n371) );
  OA22D0 U940 ( .A1(n375), .A2(n355), .B1(n376), .B2(n377), .Z(n374) );
  MUX2ND0 U941 ( .I0(n240), .I1(n154), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U942 ( .A1(n378), .A2(n373), .ZN(n240) );
  CKND2D0 U943 ( .A1(n379), .A2(n380), .ZN(n373) );
  MUX2ND0 U944 ( .I0(n380), .I1(n381), .S(n314), .ZN(n378) );
  NR2D0 U945 ( .A1(n379), .A2(n380), .ZN(n381) );
  CKND0 U946 ( .I(n382), .ZN(n379) );
  MUX2D0 U947 ( .I0(n383), .I1(n154), .S(n6), .Z(n380) );
  OA22D0 U948 ( .A1(n376), .A2(n384), .B1(n375), .B2(n359), .Z(n383) );
  MUX2ND0 U949 ( .I0(n227), .I1(n30), .S(fma_byp), .ZN(comp_mantissa_c[13]) );
  CKND2D0 U950 ( .A1(n385), .A2(n382), .ZN(n227) );
  CKND2D0 U951 ( .A1(n386), .A2(n387), .ZN(n382) );
  MUX2ND0 U952 ( .I0(n387), .I1(n388), .S(n314), .ZN(n385) );
  NR2D0 U953 ( .A1(n386), .A2(n387), .ZN(n388) );
  CKND0 U954 ( .I(n389), .ZN(n386) );
  MUX2ND0 U955 ( .I0(c[3]), .I1(n390), .S(exp_ab_greater), .ZN(n387) );
  OAI22D0 U956 ( .A1(n365), .A2(n375), .B1(n391), .B2(n376), .ZN(n390) );
  MUX2ND0 U957 ( .I0(n237), .I1(n178), .S(fma_byp), .ZN(comp_mantissa_c[12])
         );
  CKND2D0 U958 ( .A1(n392), .A2(n389), .ZN(n237) );
  CKND2D0 U959 ( .A1(n393), .A2(n394), .ZN(n389) );
  MUX2ND0 U960 ( .I0(n394), .I1(n395), .S(n314), .ZN(n392) );
  NR2D0 U961 ( .A1(n393), .A2(n394), .ZN(n395) );
  CKND0 U962 ( .I(n396), .ZN(n393) );
  OAI22D0 U963 ( .A1(exp_ab_greater), .A2(c[2]), .B1(n397), .B2(n398), .ZN(
        n394) );
  OAI32D0 U964 ( .A1(n350), .A2(n92), .A3(n399), .B1(n400), .B2(n375), .ZN(
        n398) );
  AOI21D0 U965 ( .A1(n401), .A2(exp_ab_greater), .B(n351), .ZN(n397) );
  MUX2ND0 U966 ( .I0(n228), .I1(n34), .S(fma_byp), .ZN(comp_mantissa_c[11]) );
  CKND2D0 U967 ( .A1(n402), .A2(n396), .ZN(n228) );
  CKND2D0 U968 ( .A1(n403), .A2(n404), .ZN(n396) );
  MUX2ND0 U969 ( .I0(n404), .I1(n405), .S(n314), .ZN(n402) );
  NR2D0 U970 ( .A1(n403), .A2(n404), .ZN(n405) );
  OAI21D0 U971 ( .A1(exp_ab_greater), .A2(c[1]), .B(n406), .ZN(n404) );
  OAI222D0 U972 ( .A1(n377), .A2(n375), .B1(n355), .B2(n399), .C1(n407), .C2(
        n351), .ZN(n406) );
  NR2D0 U973 ( .A1(n6), .A2(n408), .ZN(n407) );
  MUX2D0 U974 ( .I0(c[0]), .I1(n230), .S(n71), .Z(comp_mantissa_c[10]) );
  INR2D0 U975 ( .A1(n409), .B1(n403), .ZN(n230) );
  INR3D0 U976 ( .A1(n410), .B1(n906), .B2(n311), .ZN(n403) );
  CKND0 U977 ( .I(n308), .ZN(n906) );
  MUX2ND0 U978 ( .I0(n411), .I1(n2), .S(n410), .ZN(n409) );
  OAI21D0 U979 ( .A1(exp_ab_greater), .A2(c[0]), .B(n412), .ZN(n410) );
  OAI222D0 U980 ( .A1(n384), .A2(n375), .B1(n359), .B2(n399), .C1(n413), .C2(
        n351), .ZN(n412) );
  CKND0 U981 ( .I(n354), .ZN(n351) );
  CKND2D0 U982 ( .A1(exp_ab_greater), .A2(n376), .ZN(n354) );
  NR2D0 U983 ( .A1(n6), .A2(n414), .ZN(n413) );
  OAI21D0 U984 ( .A1(n2), .A2(n308), .B(n309), .ZN(n411) );
  CKND2D0 U985 ( .A1(n314), .A2(n311), .ZN(n309) );
  CKND2D0 U986 ( .A1(n315), .A2(n312), .ZN(n311) );
  CKND2D0 U987 ( .A1(exp_ab_greater), .A2(n415), .ZN(n312) );
  OAI222D0 U988 ( .A1(n416), .A2(n376), .B1(n368), .B2(n417), .C1(n401), .C2(
        n375), .ZN(n415) );
  CKND2D0 U989 ( .A1(exp_diff[3]), .A2(n418), .ZN(n417) );
  CKND0 U990 ( .I(n317), .ZN(n315) );
  CKND2D0 U991 ( .A1(n320), .A2(n318), .ZN(n317) );
  CKND2D0 U992 ( .A1(exp_ab_greater), .A2(n419), .ZN(n318) );
  OAI221D0 U993 ( .A1(n420), .A2(n375), .B1(n377), .B2(n399), .C(n421), .ZN(
        n419) );
  OA32D0 U994 ( .A1(n422), .A2(n200), .A3(n376), .B1(n423), .B2(n355), .Z(n421) );
  AOI21D0 U995 ( .A1(n325), .A2(exp_ab_greater), .B(n324), .ZN(n320) );
  CKND2D0 U996 ( .A1(n336), .A2(n424), .ZN(n324) );
  OAI21D0 U997 ( .A1(n330), .A2(n333), .B(exp_ab_greater), .ZN(n424) );
  OAI221D0 U998 ( .A1(n401), .A2(n399), .B1(n400), .B2(n423), .C(n425), .ZN(
        n333) );
  OA32D0 U999 ( .A1(n350), .A2(n92), .A3(n426), .B1(n375), .B2(n416), .Z(n425)
         );
  OAI222D0 U1000 ( .A1(n391), .A2(n399), .B1(n427), .B2(n375), .C1(n365), .C2(
        n423), .ZN(n330) );
  CKND0 U1001 ( .I(n332), .ZN(n336) );
  OAI21D0 U1002 ( .A1(n338), .A2(n6), .B(n340), .ZN(n332) );
  AOI211D0 U1003 ( .A1(n343), .A2(exp_ab_greater), .B(n532), .C(n428), .ZN(
        n340) );
  CKND0 U1004 ( .I(n298), .ZN(n428) );
  CKND0 U1005 ( .I(n344), .ZN(n532) );
  CKND2D0 U1006 ( .A1(exp_ab_greater), .A2(n429), .ZN(n344) );
  OAI222D0 U1007 ( .A1(n391), .A2(n423), .B1(n427), .B2(n399), .C1(n365), .C2(
        n426), .ZN(n429) );
  OAI222D0 U1008 ( .A1(n430), .A2(n399), .B1(n359), .B2(n426), .C1(n384), .C2(
        n423), .ZN(n343) );
  OA221D0 U1009 ( .A1(n420), .A2(n399), .B1(n377), .B2(n423), .C(n431), .Z(
        n338) );
  OA32D0 U1010 ( .A1(n422), .A2(n200), .A3(n375), .B1(n426), .B2(n355), .Z(
        n431) );
  AOI22D0 U1011 ( .A1(c[9]), .A2(n432), .B1(n433), .B2(n434), .ZN(n355) );
  ND3D0 U1012 ( .A1(n435), .A2(n436), .A3(exp_diff[4]), .ZN(n426) );
  OA221D0 U1013 ( .A1(n22), .A2(n350), .B1(n14), .B2(n422), .C(n437), .Z(n377)
         );
  AOI22D0 U1014 ( .A1(n438), .A2(c[7]), .B1(n434), .B2(c[6]), .ZN(n437) );
  CKND0 U1015 ( .I(n408), .ZN(n420) );
  OAI221D0 U1016 ( .A1(n34), .A2(n350), .B1(n154), .B2(n422), .C(n439), .ZN(
        n408) );
  AOI22D0 U1017 ( .A1(n438), .A2(c[3]), .B1(n434), .B2(c[2]), .ZN(n439) );
  CKND0 U1018 ( .I(c[1]), .ZN(n34) );
  OAI222D0 U1019 ( .A1(n359), .A2(n423), .B1(n430), .B2(n375), .C1(n384), .C2(
        n399), .ZN(n325) );
  OA221D0 U1020 ( .A1(n154), .A2(n350), .B1(n124), .B2(n422), .C(n440), .Z(
        n384) );
  AOI22D0 U1021 ( .A1(n438), .A2(c[6]), .B1(n434), .B2(c[5]), .ZN(n440) );
  CKND0 U1022 ( .I(c[4]), .ZN(n154) );
  CKND0 U1023 ( .I(n414), .ZN(n430) );
  OAI221D0 U1024 ( .A1(n200), .A2(n350), .B1(n30), .B2(n422), .C(n441), .ZN(
        n414) );
  AOI22D0 U1025 ( .A1(n438), .A2(c[2]), .B1(n434), .B2(c[1]), .ZN(n441) );
  CKND0 U1026 ( .I(c[3]), .ZN(n30) );
  CKND0 U1027 ( .I(c[0]), .ZN(n200) );
  AOI222D0 U1028 ( .A1(c[8]), .A2(n432), .B1(n433), .B2(n438), .C1(c[9]), .C2(
        n434), .ZN(n359) );
  CKND0 U1029 ( .I(n2), .ZN(n314) );
  CKND2D0 U1030 ( .A1(exp_ab_greater), .A2(n442), .ZN(n308) );
  OAI222D0 U1031 ( .A1(n391), .A2(n375), .B1(n427), .B2(n376), .C1(n365), .C2(
        n399), .ZN(n442) );
  OA221D0 U1032 ( .A1(n92), .A2(n422), .B1(n124), .B2(n350), .C(n443), .Z(n365) );
  AOI22D0 U1033 ( .A1(n434), .A2(c[8]), .B1(n438), .B2(c[9]), .ZN(n443) );
  CKND0 U1034 ( .I(c[7]), .ZN(n124) );
  CKND0 U1035 ( .I(n433), .ZN(n92) );
  ND3D0 U1036 ( .A1(n436), .A2(n418), .A3(n435), .ZN(n376) );
  AOI222D0 U1037 ( .A1(c[2]), .A2(n444), .B1(n434), .B2(c[0]), .C1(c[1]), .C2(
        n438), .ZN(n427) );
  ND3D0 U1038 ( .A1(n436), .A2(n418), .A3(exp_diff[2]), .ZN(n375) );
  OA221D0 U1039 ( .A1(n23), .A2(n422), .B1(n22), .B2(n445), .C(n446), .Z(n391)
         );
  AOI22D0 U1040 ( .A1(n432), .A2(c[3]), .B1(n434), .B2(c[4]), .ZN(n446) );
  CKND0 U1041 ( .I(c[6]), .ZN(n23) );
  CKND2D0 U1042 ( .A1(c[15]), .A2(n5), .ZN(n2) );
  CKND0 U1043 ( .I(add_byp), .ZN(n5) );
  NR2D0 U1044 ( .A1(fma_byp), .A2(n298), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n447), .ZN(n298) );
  OAI222D0 U1046 ( .A1(n416), .A2(n399), .B1(n368), .B2(n448), .C1(n401), .C2(
        n423), .ZN(n447) );
  ND3D0 U1047 ( .A1(exp_diff[3]), .A2(n418), .A3(exp_diff[2]), .ZN(n423) );
  OA221D0 U1048 ( .A1(n178), .A2(n350), .B1(n22), .B2(n422), .C(n449), .Z(n401) );
  AOI22D0 U1049 ( .A1(n438), .A2(c[4]), .B1(n434), .B2(c[3]), .ZN(n449) );
  CKND0 U1050 ( .I(c[5]), .ZN(n22) );
  CKND0 U1051 ( .I(n432), .ZN(n350) );
  CKND0 U1052 ( .I(c[2]), .ZN(n178) );
  CKND2D0 U1053 ( .A1(exp_diff[4]), .A2(n436), .ZN(n448) );
  CKND0 U1054 ( .I(exp_diff[3]), .ZN(n436) );
  MUX2D0 U1055 ( .I0(n450), .I1(n400), .S(n435), .Z(n368) );
  OA221D0 U1056 ( .A1(n15), .A2(n422), .B1(n14), .B2(n445), .C(n451), .Z(n400)
         );
  AOI22D0 U1057 ( .A1(n432), .A2(c[6]), .B1(n434), .B2(c[7]), .ZN(n451) );
  NR2D0 U1058 ( .A1(n452), .A2(exp_diff[1]), .ZN(n434) );
  CKND0 U1059 ( .I(c[8]), .ZN(n14) );
  CKND0 U1060 ( .I(c[9]), .ZN(n15) );
  CKND2D0 U1061 ( .A1(n432), .A2(n433), .ZN(n450) );
  ND4D0 U1062 ( .A1(n305), .A2(n303), .A3(n453), .A4(n301), .ZN(n433) );
  CKND0 U1063 ( .I(c[12]), .ZN(n301) );
  NR2D0 U1064 ( .A1(c[14]), .A2(c[13]), .ZN(n453) );
  CKND0 U1065 ( .I(c[11]), .ZN(n303) );
  CKND0 U1066 ( .I(c[10]), .ZN(n305) );
  NR2D0 U1067 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n432) );
  ND3D0 U1068 ( .A1(n435), .A2(n418), .A3(exp_diff[3]), .ZN(n399) );
  CKND0 U1069 ( .I(exp_diff[4]), .ZN(n418) );
  CKND0 U1070 ( .I(exp_diff[2]), .ZN(n435) );
  AOI22D0 U1071 ( .A1(c[1]), .A2(n444), .B1(c[0]), .B2(n438), .ZN(n416) );
  CKND0 U1072 ( .I(n445), .ZN(n438) );
  CKND2D0 U1073 ( .A1(exp_diff[1]), .A2(n452), .ZN(n445) );
  CKND0 U1074 ( .I(exp_diff[0]), .ZN(n452) );
  CKND0 U1075 ( .I(n422), .ZN(n444) );
  CKND2D0 U1076 ( .A1(exp_diff[1]), .A2(exp_diff[0]), .ZN(n422) );
  MUX2ND0 U1077 ( .I0(n231), .I1(n13), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1078 ( .I(mantissa_ab[9]), .ZN(n13) );
  CKXOR2D0 U1079 ( .A1(n1063), .A2(n454), .Z(n231) );
  CKND0 U1080 ( .I(n455), .ZN(n1063) );
  MUX2D0 U1081 ( .I0(mantissa_ab[8]), .I1(n244), .S(n71), .Z(
        comp_mantissa_ab[8]) );
  AN2D0 U1082 ( .A1(n456), .A2(n457), .Z(n244) );
  MUX2ND0 U1083 ( .I0(n458), .I1(n459), .S(sign_ab), .ZN(n456) );
  NR2D0 U1084 ( .A1(n460), .A2(n458), .ZN(n459) );
  MUX2ND0 U1085 ( .I0(n245), .I1(n19), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1086 ( .I(mantissa_ab[7]), .ZN(n19) );
  CKND2D0 U1087 ( .A1(n461), .A2(n462), .ZN(n245) );
  MUX2ND0 U1088 ( .I0(n463), .I1(n464), .S(sign_ab), .ZN(n461) );
  NR2D0 U1089 ( .A1(n465), .A2(n463), .ZN(n464) );
  MUX2ND0 U1090 ( .I0(n255), .I1(n20), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1091 ( .I(mantissa_ab[6]), .ZN(n20) );
  CKND2D0 U1092 ( .A1(n466), .A2(n467), .ZN(n255) );
  MUX2ND0 U1093 ( .I0(n468), .I1(n469), .S(sign_ab), .ZN(n466) );
  NR2D0 U1094 ( .A1(n470), .A2(n468), .ZN(n469) );
  MUX2ND0 U1095 ( .I0(n282), .I1(n37), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1096 ( .I(mantissa_ab[5]), .ZN(n37) );
  CKND2D0 U1097 ( .A1(n471), .A2(n472), .ZN(n282) );
  MUX2ND0 U1098 ( .I0(n473), .I1(n474), .S(sign_ab), .ZN(n471) );
  NR2D0 U1099 ( .A1(n475), .A2(n473), .ZN(n474) );
  MUX2ND0 U1100 ( .I0(n285), .I1(n26), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1101 ( .I(mantissa_ab[4]), .ZN(n26) );
  CKND2D0 U1102 ( .A1(n476), .A2(n477), .ZN(n285) );
  MUX2ND0 U1103 ( .I0(n478), .I1(n479), .S(sign_ab), .ZN(n476) );
  NR2D0 U1104 ( .A1(n480), .A2(n478), .ZN(n479) );
  MUX2D0 U1105 ( .I0(mantissa_ab[3]), .I1(n274), .S(n71), .Z(
        comp_mantissa_ab[3]) );
  INR2D0 U1106 ( .A1(n481), .B1(n480), .ZN(n274) );
  MUX2ND0 U1107 ( .I0(n482), .I1(n483), .S(sign_ab), .ZN(n481) );
  NR2D0 U1108 ( .A1(n484), .A2(n482), .ZN(n483) );
  MUX2D0 U1109 ( .I0(mantissa_ab[2]), .I1(n267), .S(n71), .Z(
        comp_mantissa_ab[2]) );
  INR2D0 U1110 ( .A1(n485), .B1(n484), .ZN(n267) );
  MUX2ND0 U1111 ( .I0(n486), .I1(n8), .S(n487), .ZN(n485) );
  NR2D0 U1112 ( .A1(n209), .A2(fma_byp), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1113 ( .A1(n488), .A2(n530), .A3(n531), .B(sign_ab), .ZN(n209) );
  CKND0 U1114 ( .I(n489), .ZN(n530) );
  MUX2ND0 U1115 ( .I0(n96), .I1(n490), .S(fma_byp), .ZN(comp_mantissa_ab[20])
         );
  CKND0 U1116 ( .I(N800), .ZN(n490) );
  XNR2D0 U1117 ( .A1(n1103), .A2(n531), .ZN(n96) );
  MUX2D0 U1118 ( .I0(N800), .I1(N65), .S(n307), .Z(n531) );
  OAI21D0 U1119 ( .A1(n8), .A2(n489), .B(n491), .ZN(n1103) );
  MUX2ND0 U1120 ( .I0(n271), .I1(n492), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1121 ( .I(mantissa_ab[1]), .ZN(n492) );
  MUX2ND0 U1122 ( .I0(n493), .I1(n486), .S(n296), .ZN(n271) );
  CKND0 U1123 ( .I(n295), .ZN(n486) );
  CKND2D0 U1124 ( .A1(sign_ab), .A2(n494), .ZN(n295) );
  IND2D0 U1125 ( .A1(n297), .B1(sign_ab), .ZN(n493) );
  MUX2ND0 U1126 ( .I0(n108), .I1(n495), .S(fma_byp), .ZN(comp_mantissa_ab[19])
         );
  CKND0 U1127 ( .I(mantissa_ab[19]), .ZN(n495) );
  CKXOR2D0 U1128 ( .A1(n529), .A2(n489), .Z(n108) );
  MUX2ND0 U1129 ( .I0(mantissa_ab[19]), .I1(N64), .S(n307), .ZN(n489) );
  CKND0 U1130 ( .I(n491), .ZN(n529) );
  CKND2D0 U1131 ( .A1(sign_ab), .A2(n488), .ZN(n491) );
  ND3D0 U1132 ( .A1(n496), .A2(n497), .A3(n498), .ZN(n488) );
  MUX2D0 U1133 ( .I0(mantissa_ab[18]), .I1(n116), .S(n71), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1134 ( .A1(n499), .A2(n497), .ZN(n116) );
  MUX2ND0 U1135 ( .I0(mantissa_ab[18]), .I1(N63), .S(n307), .ZN(n497) );
  AOI21D0 U1136 ( .A1(n498), .A2(n496), .B(n8), .ZN(n499) );
  MUX2D0 U1137 ( .I0(mantissa_ab[17]), .I1(n129), .S(n71), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1138 ( .A1(n500), .A2(n496), .ZN(n129) );
  MUX2ND0 U1139 ( .I0(mantissa_ab[17]), .I1(N62), .S(n307), .ZN(n496) );
  NR2D0 U1140 ( .A1(n498), .A2(n8), .ZN(n500) );
  INR2D0 U1141 ( .A1(n501), .B1(n502), .ZN(n498) );
  MUX2D0 U1142 ( .I0(mantissa_ab[16]), .I1(n138), .S(n71), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1143 ( .A1(n503), .A2(n501), .ZN(n138) );
  MUX2ND0 U1144 ( .I0(mantissa_ab[16]), .I1(N61), .S(n307), .ZN(n501) );
  INR2D0 U1145 ( .A1(n502), .B1(n8), .ZN(n503) );
  MUX2ND0 U1146 ( .I0(n148), .I1(n504), .S(fma_byp), .ZN(comp_mantissa_ab[15])
         );
  CKND0 U1147 ( .I(mantissa_ab[15]), .ZN(n504) );
  CKND2D0 U1148 ( .A1(n505), .A2(n502), .ZN(n148) );
  CKND2D0 U1149 ( .A1(n506), .A2(n507), .ZN(n502) );
  MUX2ND0 U1150 ( .I0(n507), .I1(n508), .S(sign_ab), .ZN(n505) );
  NR2D0 U1151 ( .A1(n506), .A2(n507), .ZN(n508) );
  CKND0 U1152 ( .I(n509), .ZN(n506) );
  MUX2ND0 U1153 ( .I0(N60), .I1(mantissa_ab[15]), .S(n12), .ZN(n507) );
  MUX2D0 U1154 ( .I0(mantissa_ab[14]), .I1(n238), .S(n71), .Z(
        comp_mantissa_ab[14]) );
  CKND0 U1155 ( .I(n158), .ZN(n238) );
  CKND2D0 U1156 ( .A1(n510), .A2(n509), .ZN(n158) );
  CKND2D0 U1157 ( .A1(n511), .A2(n512), .ZN(n509) );
  MUX2ND0 U1158 ( .I0(n512), .I1(n513), .S(sign_ab), .ZN(n510) );
  NR2D0 U1159 ( .A1(n511), .A2(n512), .ZN(n513) );
  AN2D0 U1160 ( .A1(n514), .A2(n515), .Z(n511) );
  MUX2ND0 U1161 ( .I0(N59), .I1(mantissa_ab[14]), .S(n12), .ZN(n512) );
  MUX2D0 U1162 ( .I0(mantissa_ab[13]), .I1(n173), .S(n71), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1163 ( .A1(n516), .A2(n515), .ZN(n173) );
  MUX2ND0 U1164 ( .I0(mantissa_ab[13]), .I1(N58), .S(n307), .ZN(n515) );
  NR2D0 U1165 ( .A1(n514), .A2(n8), .ZN(n516) );
  INR2D0 U1166 ( .A1(n517), .B1(n518), .ZN(n514) );
  MUX2D0 U1167 ( .I0(mantissa_ab[12]), .I1(n183), .S(n71), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1168 ( .A1(n519), .A2(n517), .ZN(n183) );
  MUX2ND0 U1169 ( .I0(mantissa_ab[12]), .I1(N57), .S(n307), .ZN(n517) );
  INR2D0 U1170 ( .A1(n518), .B1(n8), .ZN(n519) );
  MUX2ND0 U1171 ( .I0(n192), .I1(n520), .S(fma_byp), .ZN(comp_mantissa_ab[11])
         );
  CKND0 U1172 ( .I(mantissa_ab[11]), .ZN(n520) );
  CKND2D0 U1173 ( .A1(n521), .A2(n518), .ZN(n192) );
  CKND2D0 U1174 ( .A1(n522), .A2(n523), .ZN(n518) );
  MUX2ND0 U1175 ( .I0(n523), .I1(n524), .S(sign_ab), .ZN(n521) );
  NR2D0 U1176 ( .A1(n522), .A2(n523), .ZN(n524) );
  MUX2ND0 U1177 ( .I0(N56), .I1(mantissa_ab[11]), .S(n12), .ZN(n523) );
  MUX2D0 U1178 ( .I0(mantissa_ab[10]), .I1(n205), .S(n71), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1179 ( .I(fma_byp), .ZN(n71) );
  INR2D0 U1180 ( .A1(n525), .B1(n522), .ZN(n205) );
  INR3D0 U1181 ( .A1(n526), .B1(n544), .B2(n457), .ZN(n522) );
  CKND0 U1182 ( .I(n454), .ZN(n544) );
  MUX2ND0 U1183 ( .I0(n527), .I1(n8), .S(n526), .ZN(n525) );
  MUX2ND0 U1184 ( .I0(N55), .I1(mantissa_ab[10]), .S(n12), .ZN(n526) );
  OAI21D0 U1185 ( .A1(n454), .A2(n8), .B(n455), .ZN(n527) );
  CKND2D0 U1186 ( .A1(sign_ab), .A2(n457), .ZN(n455) );
  CKND2D0 U1187 ( .A1(n460), .A2(n458), .ZN(n457) );
  MUX2ND0 U1188 ( .I0(N53), .I1(mantissa_ab[8]), .S(n12), .ZN(n458) );
  CKND0 U1189 ( .I(n462), .ZN(n460) );
  CKND2D0 U1190 ( .A1(n465), .A2(n463), .ZN(n462) );
  MUX2ND0 U1191 ( .I0(N52), .I1(mantissa_ab[7]), .S(n12), .ZN(n463) );
  CKND0 U1192 ( .I(n467), .ZN(n465) );
  CKND2D0 U1193 ( .A1(n470), .A2(n468), .ZN(n467) );
  MUX2ND0 U1194 ( .I0(N51), .I1(mantissa_ab[6]), .S(n12), .ZN(n468) );
  CKND0 U1195 ( .I(n472), .ZN(n470) );
  CKND2D0 U1196 ( .A1(n475), .A2(n473), .ZN(n472) );
  MUX2ND0 U1197 ( .I0(N50), .I1(mantissa_ab[5]), .S(n12), .ZN(n473) );
  CKND0 U1198 ( .I(n477), .ZN(n475) );
  CKND2D0 U1199 ( .A1(n480), .A2(n478), .ZN(n477) );
  MUX2ND0 U1200 ( .I0(N49), .I1(mantissa_ab[4]), .S(n12), .ZN(n478) );
  AN2D0 U1201 ( .A1(n484), .A2(n482), .Z(n480) );
  MUX2ND0 U1202 ( .I0(N48), .I1(mantissa_ab[3]), .S(n12), .ZN(n482) );
  INR2D0 U1203 ( .A1(n487), .B1(n494), .ZN(n484) );
  CKND2D0 U1218 ( .A1(n297), .A2(n296), .ZN(n494) );
  MUX2ND0 U1219 ( .I0(N46), .I1(mantissa_ab[1]), .S(n12), .ZN(n296) );
  MUX2ND0 U1220 ( .I0(N47), .I1(mantissa_ab[2]), .S(n12), .ZN(n487) );
  CKND0 U1221 ( .I(sign_ab), .ZN(n8) );
  MUX2ND0 U1222 ( .I0(mantissa_ab[9]), .I1(N54), .S(n307), .ZN(n454) );
  MUX2ND0 U1223 ( .I0(n297), .I1(n36), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1224 ( .I(mantissa_ab[0]), .ZN(n36) );
  MUX2ND0 U1225 ( .I0(mantissa_ab[0]), .I1(N45), .S(n307), .ZN(n297) );
  CKND0 U1226 ( .I(n12), .ZN(n307) );
  CKND2D0 U1227 ( .A1(exp_ab_less), .A2(n6), .ZN(n12) );
  CKND0 U1228 ( .I(exp_ab_greater), .ZN(n6) );
  ND4D0 U1229 ( .A1(n306), .A2(n304), .A3(n528), .A4(n302), .ZN(N800) );
  CKND0 U1230 ( .I(exp_ab[2]), .ZN(n302) );
  NR2D0 U1231 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n528) );
  CKND0 U1232 ( .I(exp_ab[1]), .ZN(n304) );
  CKND0 U1233 ( .I(exp_ab[0]), .ZN(n306) );
endmodule


module fma_normalizer_rounder_1_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [19:0] A;
  input [4:0] SH;
  output [19:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][3] ,
         \ML_int[4][2] , \ML_int[4][1] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2D0 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2D0 M1_1_18 ( .I0(\ML_int[1][18] ), .I1(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2D0 M1_2_18 ( .I0(\ML_int[2][18] ), .I1(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2D0 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2D0 M1_1_19 ( .I0(\ML_int[1][19] ), .I1(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2D0 M1_2_19 ( .I0(\ML_int[2][19] ), .I1(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2D0 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2D0 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2D0 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2D0 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2D0 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2D0 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2D0 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2D0 M1_3_19 ( .I0(\ML_int[3][19] ), .I1(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2D0 M1_4_19 ( .I0(\ML_int[4][19] ), .I1(\ML_int[4][3] ), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2D0 M1_3_18 ( .I0(\ML_int[3][18] ), .I1(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2D0 M1_4_18 ( .I0(\ML_int[4][18] ), .I1(\ML_int[4][2] ), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2D0 M1_3_17 ( .I0(\ML_int[3][17] ), .I1(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2D0 M1_4_17 ( .I0(\ML_int[4][17] ), .I1(\ML_int[4][1] ), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2D0 M1_1_16 ( .I0(\ML_int[1][16] ), .I1(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2D0 M1_2_16 ( .I0(\ML_int[2][16] ), .I1(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2D0 M1_1_17 ( .I0(\ML_int[1][17] ), .I1(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2D0 M1_2_17 ( .I0(\ML_int[2][17] ), .I1(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2D0 M1_2_4 ( .I0(\ML_int[2][4] ), .I1(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2D0 M1_2_5 ( .I0(\ML_int[2][5] ), .I1(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0 M1_2_6 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2D0 M1_2_7 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2D0 M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D0 M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2D0 M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D0 M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2D0 M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0 M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0 M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2D0 M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0 M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2D0 M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0 M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0 M1_1_13 ( .I0(\ML_int[1][13] ), .I1(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2D0 M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0 M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0 M1_1_14 ( .I0(\ML_int[1][14] ), .I1(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2D0 M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2D0 M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0 M1_1_15 ( .I0(\ML_int[1][15] ), .I1(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2D0 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0 M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2D0 M1_2_13 ( .I0(\ML_int[2][13] ), .I1(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2D0 M1_2_14 ( .I0(\ML_int[2][14] ), .I1(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2D0 M1_2_15 ( .I0(\ML_int[2][15] ), .I1(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  INVD1 U3 ( .I(n18), .ZN(n9) );
  INVD1 U4 ( .I(n16), .ZN(n10) );
  INVD1 U5 ( .I(n17), .ZN(n11) );
  INVD1 U6 ( .I(SH[3]), .ZN(n14) );
  INVD1 U7 ( .I(SH[2]), .ZN(n12) );
  INVD1 U8 ( .I(SH[1]), .ZN(n13) );
  NR2D1 U9 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][9] ) );
  MUX2ND0 U10 ( .I0(\ML_int[3][9] ), .I1(n9), .S(SH[3]), .ZN(n1) );
  NR2D1 U11 ( .A1(n2), .A2(SH[4]), .ZN(\ML_int[5][14] ) );
  MUX2ND0 U12 ( .I0(\ML_int[3][14] ), .I1(\ML_int[3][6] ), .S(SH[3]), .ZN(n2)
         );
  NR2D1 U13 ( .A1(n3), .A2(SH[4]), .ZN(\ML_int[5][10] ) );
  MUX2ND0 U14 ( .I0(\ML_int[3][10] ), .I1(n11), .S(SH[3]), .ZN(n3) );
  NR2D1 U15 ( .A1(n4), .A2(SH[4]), .ZN(\ML_int[5][15] ) );
  MUX2ND0 U16 ( .I0(\ML_int[3][15] ), .I1(\ML_int[3][7] ), .S(SH[3]), .ZN(n4)
         );
  NR2D1 U17 ( .A1(n5), .A2(SH[4]), .ZN(\ML_int[5][12] ) );
  MUX2ND0 U18 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), .ZN(n5)
         );
  NR2D1 U19 ( .A1(n6), .A2(SH[4]), .ZN(\ML_int[5][11] ) );
  MUX2ND0 U20 ( .I0(\ML_int[3][11] ), .I1(n10), .S(SH[3]), .ZN(n6) );
  MUX2ND0 U21 ( .I0(n7), .I1(n15), .S(SH[4]), .ZN(\ML_int[5][16] ) );
  MUX2ND0 U22 ( .I0(\ML_int[3][16] ), .I1(\ML_int[3][8] ), .S(SH[3]), .ZN(n7)
         );
  NR2D1 U23 ( .A1(n8), .A2(SH[4]), .ZN(\ML_int[5][13] ) );
  MUX2ND0 U24 ( .I0(\ML_int[3][13] ), .I1(\ML_int[3][5] ), .S(SH[3]), .ZN(n8)
         );
  INR2D1 U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  NR2D0 U26 ( .A1(SH[4]), .A2(n15), .ZN(\ML_int[5][0] ) );
  NR2D0 U27 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][3] ) );
  NR2D0 U28 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][2] ) );
  NR2D0 U29 ( .A1(SH[3]), .A2(n18), .ZN(\ML_int[4][1] ) );
  ND3D0 U30 ( .A1(n12), .A2(n14), .A3(\ML_int[2][0] ), .ZN(n15) );
  CKND2D0 U31 ( .A1(\ML_int[2][3] ), .A2(n12), .ZN(n16) );
  CKND2D0 U32 ( .A1(\ML_int[2][2] ), .A2(n12), .ZN(n17) );
  CKND2D0 U33 ( .A1(\ML_int[2][1] ), .A2(n12), .ZN(n18) );
  AN2D0 U34 ( .A1(\ML_int[1][1] ), .A2(n13), .Z(\ML_int[2][1] ) );
  AN2D0 U35 ( .A1(\ML_int[1][0] ), .A2(n13), .Z(\ML_int[2][0] ) );
endmodule


module fma_normalizer_rounder_1_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1 U1_4 ( .A1(A[4]), .A2(B_AS[4]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1D0 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1D0 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1D0 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0])
         );
  CKXOR2D0 U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0 U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0 U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0 U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0 U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module fma_normalizer_rounder_1 ( mantissa_ab_c_in, exp_ab_c_in, 
        mantissa_shift, fma_byp, rounder_start, mantissa_ab_c_out, 
        exp_ab_c_out, rounder_done );
  input [21:0] mantissa_ab_c_in;
  input [4:0] exp_ab_c_in;
  input [4:0] mantissa_shift;
  output [9:0] mantissa_ab_c_out;
  output [4:0] exp_ab_c_out;
  input fma_byp, rounder_start;
  output rounder_done;
  wire   rounder_start, N11, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign rounder_done = rounder_start;

  fma_normalizer_rounder_1_DW01_ash_0 sll_926 ( .A(mantissa_ab_c_in[19:0]), 
        .DATA_TC(n78), .SH({n77, n76, n74, n75, N11}), .SH_TC(n78), .B({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N24}) );
  fma_normalizer_rounder_1_DW01_addsub_0 r82 ( .A(exp_ab_c_in), .B({
        \U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), 
        .CI(n78), .ADD_SUB(\U3/U2/Z_0 ), .SUM({N23, N22, N21, N20, N19}) );
  TIEL U3 ( .ZN(n78) );
  CKND0 U4 ( .I(n1), .ZN(n74) );
  CKND0 U5 ( .I(n2), .ZN(n75) );
  CKND0 U6 ( .I(n3), .ZN(n76) );
  CKND0 U7 ( .I(n4), .ZN(n77) );
  IOA21D0 U8 ( .A1(fma_byp), .A2(mantissa_ab_c_in[19]), .B(n5), .ZN(
        mantissa_ab_c_out[9]) );
  MUX2ND0 U9 ( .I0(n6), .I1(n7), .S(n8), .ZN(n5) );
  OAI21D0 U10 ( .A1(n9), .A2(n10), .B(n11), .ZN(n7) );
  AN2D0 U11 ( .A1(n10), .A2(n12), .Z(n6) );
  IOA21D0 U12 ( .A1(fma_byp), .A2(mantissa_ab_c_in[18]), .B(n13), .ZN(
        mantissa_ab_c_out[8]) );
  MUX2ND0 U13 ( .I0(n12), .I1(n14), .S(n10), .ZN(n13) );
  CKND0 U14 ( .I(n11), .ZN(n14) );
  AOI21D0 U15 ( .A1(n15), .A2(n16), .B(n17), .ZN(n11) );
  IOA21D0 U16 ( .A1(fma_byp), .A2(mantissa_ab_c_in[17]), .B(n18), .ZN(
        mantissa_ab_c_out[7]) );
  MUX2ND0 U17 ( .I0(n17), .I1(n19), .S(n16), .ZN(n18) );
  NR2D0 U18 ( .A1(n9), .A2(n20), .ZN(n19) );
  OAI21D0 U19 ( .A1(n21), .A2(n9), .B(n22), .ZN(n17) );
  IOA21D0 U20 ( .A1(fma_byp), .A2(mantissa_ab_c_in[16]), .B(n24), .ZN(
        mantissa_ab_c_out[6]) );
  MUX2ND0 U21 ( .I0(n25), .I1(n26), .S(n27), .ZN(n24) );
  NR3D0 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n26) );
  AO21D0 U23 ( .A1(n15), .A2(n30), .B(n31), .Z(n25) );
  IOA21D0 U24 ( .A1(fma_byp), .A2(mantissa_ab_c_in[15]), .B(n32), .ZN(
        mantissa_ab_c_out[5]) );
  MUX2ND0 U25 ( .I0(n31), .I1(n33), .S(n30), .ZN(n32) );
  NR2D0 U26 ( .A1(n29), .A2(n28), .ZN(n33) );
  AO21D0 U27 ( .A1(n15), .A2(n29), .B(n34), .Z(n31) );
  IOA21D0 U28 ( .A1(fma_byp), .A2(mantissa_ab_c_in[14]), .B(n35), .ZN(
        mantissa_ab_c_out[4]) );
  MUX2ND0 U29 ( .I0(n34), .I1(n36), .S(n29), .ZN(n35) );
  CKND0 U30 ( .I(n28), .ZN(n36) );
  CKND2D0 U31 ( .A1(n15), .A2(n37), .ZN(n28) );
  OAI21D0 U32 ( .A1(n37), .A2(n9), .B(n22), .ZN(n34) );
  IOA21D0 U33 ( .A1(fma_byp), .A2(mantissa_ab_c_in[13]), .B(n38), .ZN(
        mantissa_ab_c_out[3]) );
  MUX2ND0 U34 ( .I0(n39), .I1(n40), .S(n41), .ZN(n38) );
  NR3D0 U35 ( .A1(n9), .A2(n42), .A3(n43), .ZN(n40) );
  AO21D0 U36 ( .A1(n15), .A2(n42), .B(n44), .Z(n39) );
  IOA21D0 U37 ( .A1(fma_byp), .A2(mantissa_ab_c_in[12]), .B(n45), .ZN(
        mantissa_ab_c_out[2]) );
  MUX2ND0 U38 ( .I0(n44), .I1(n46), .S(n42), .ZN(n45) );
  NR2D0 U39 ( .A1(n43), .A2(n9), .ZN(n46) );
  AO21D0 U40 ( .A1(n15), .A2(n47), .B(n48), .Z(n44) );
  IOA21D0 U41 ( .A1(fma_byp), .A2(mantissa_ab_c_in[11]), .B(n49), .ZN(
        mantissa_ab_c_out[1]) );
  MUX2ND0 U42 ( .I0(n48), .I1(n50), .S(n47), .ZN(n49) );
  NR2D0 U43 ( .A1(n51), .A2(n9), .ZN(n50) );
  IOA21D0 U44 ( .A1(n51), .A2(n15), .B(n22), .ZN(n48) );
  CKND0 U45 ( .I(n52), .ZN(n22) );
  IOA21D0 U46 ( .A1(fma_byp), .A2(mantissa_ab_c_in[10]), .B(n53), .ZN(
        mantissa_ab_c_out[0]) );
  MUX2ND0 U47 ( .I0(n52), .I1(n15), .S(n51), .ZN(n53) );
  NR2D0 U48 ( .A1(n54), .A2(fma_byp), .ZN(n52) );
  MUX2ND0 U49 ( .I0(n55), .I1(n56), .S(n57), .ZN(exp_ab_c_out[4]) );
  XNR2D0 U50 ( .A1(N23), .A2(n58), .ZN(n56) );
  XNR2D0 U51 ( .A1(n58), .A2(exp_ab_c_in[4]), .ZN(n55) );
  INR3D0 U52 ( .A1(n59), .B1(n60), .B2(n61), .ZN(n58) );
  CKXOR2D0 U53 ( .A1(n62), .A2(n59), .Z(exp_ab_c_out[3]) );
  MUX2D0 U54 ( .I0(exp_ab_c_in[3]), .I1(N22), .S(n57), .Z(n59) );
  NR2D0 U55 ( .A1(n61), .A2(n60), .ZN(n62) );
  CKXOR2D0 U56 ( .A1(n60), .A2(n61), .Z(exp_ab_c_out[2]) );
  MUX2ND0 U57 ( .I0(exp_ab_c_in[2]), .I1(N21), .S(n57), .ZN(n61) );
  IND3D0 U58 ( .A1(n63), .B1(n64), .B2(n65), .ZN(n60) );
  CKXOR2D0 U59 ( .A1(n63), .A2(n66), .Z(exp_ab_c_out[1]) );
  CKND2D0 U60 ( .A1(n65), .A2(n64), .ZN(n66) );
  MUX2ND0 U61 ( .I0(exp_ab_c_in[1]), .I1(N20), .S(n57), .ZN(n63) );
  CKXOR2D0 U62 ( .A1(n65), .A2(n64), .Z(exp_ab_c_out[0]) );
  MUX2D0 U63 ( .I0(exp_ab_c_in[0]), .I1(N19), .S(n57), .Z(n64) );
  NR2D0 U64 ( .A1(n67), .A2(fma_byp), .ZN(n57) );
  AN3D0 U65 ( .A1(n8), .A2(n10), .A3(n12), .Z(n65) );
  NR3D0 U66 ( .A1(n9), .A2(n16), .A3(n20), .ZN(n12) );
  CKND0 U67 ( .I(n21), .ZN(n20) );
  INR4D0 U68 ( .A1(n37), .B1(n27), .B2(n30), .B3(n29), .ZN(n21) );
  AOI222D0 U69 ( .A1(mantissa_ab_c_in[14]), .A2(n67), .B1(mantissa_ab_c_in[15]), .B2(mantissa_ab_c_in[21]), .C1(N30), .C2(\U3/U2/Z_0 ), .ZN(n29) );
  AOI222D0 U70 ( .A1(mantissa_ab_c_in[15]), .A2(n67), .B1(mantissa_ab_c_in[16]), .B2(mantissa_ab_c_in[21]), .C1(N31), .C2(\U3/U2/Z_0 ), .ZN(n30) );
  AOI222D0 U71 ( .A1(mantissa_ab_c_in[16]), .A2(n67), .B1(mantissa_ab_c_in[17]), .B2(mantissa_ab_c_in[21]), .C1(N32), .C2(\U3/U2/Z_0 ), .ZN(n27) );
  NR3D0 U72 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n37) );
  OR2D0 U73 ( .A1(n47), .A2(n51), .Z(n43) );
  AOI222D0 U74 ( .A1(mantissa_ab_c_in[11]), .A2(n67), .B1(mantissa_ab_c_in[12]), .B2(mantissa_ab_c_in[21]), .C1(N27), .C2(\U3/U2/Z_0 ), .ZN(n47) );
  AOI222D0 U75 ( .A1(mantissa_ab_c_in[12]), .A2(n67), .B1(mantissa_ab_c_in[13]), .B2(mantissa_ab_c_in[21]), .C1(N28), .C2(\U3/U2/Z_0 ), .ZN(n42) );
  AOI222D0 U76 ( .A1(mantissa_ab_c_in[13]), .A2(n67), .B1(mantissa_ab_c_in[14]), .B2(mantissa_ab_c_in[21]), .C1(N29), .C2(\U3/U2/Z_0 ), .ZN(n41) );
  AOI222D0 U77 ( .A1(mantissa_ab_c_in[17]), .A2(n67), .B1(mantissa_ab_c_in[18]), .B2(mantissa_ab_c_in[21]), .C1(N33), .C2(\U3/U2/Z_0 ), .ZN(n16) );
  CKND0 U78 ( .I(n15), .ZN(n9) );
  INR2D0 U79 ( .A1(n54), .B1(fma_byp), .ZN(n15) );
  AOI31D0 U80 ( .A1(n51), .A2(n68), .A3(n69), .B(n70), .ZN(n54) );
  AOI222D0 U81 ( .A1(N25), .A2(\U3/U2/Z_0 ), .B1(mantissa_ab_c_in[9]), .B2(n67), .C1(mantissa_ab_c_in[10]), .C2(mantissa_ab_c_in[21]), .ZN(n70) );
  AOI22D0 U82 ( .A1(mantissa_ab_c_in[0]), .A2(n67), .B1(N24), .B2(\U3/U2/Z_0 ), 
        .ZN(n69) );
  CKND2D0 U83 ( .A1(mantissa_ab_c_in[1]), .A2(mantissa_ab_c_in[21]), .ZN(n68)
         );
  AOI222D0 U84 ( .A1(mantissa_ab_c_in[10]), .A2(n67), .B1(mantissa_ab_c_in[11]), .B2(mantissa_ab_c_in[21]), .C1(N26), .C2(\U3/U2/Z_0 ), .ZN(n51) );
  AO222D0 U85 ( .A1(mantissa_ab_c_in[18]), .A2(n67), .B1(mantissa_ab_c_in[21]), 
        .B2(mantissa_ab_c_in[19]), .C1(N34), .C2(\U3/U2/Z_0 ), .Z(n10) );
  AO222D0 U86 ( .A1(n67), .A2(mantissa_ab_c_in[19]), .B1(mantissa_ab_c_in[20]), 
        .B2(mantissa_ab_c_in[21]), .C1(N35), .C2(\U3/U2/Z_0 ), .Z(n8) );
  NR2D0 U87 ( .A1(\U3/U2/Z_0 ), .A2(mantissa_ab_c_in[21]), .ZN(n67) );
  NR2D0 U88 ( .A1(n71), .A2(n4), .ZN(\U3/U1/Z_4 ) );
  CKND2D0 U89 ( .A1(mantissa_shift[4]), .A2(n72), .ZN(n4) );
  NR2D0 U90 ( .A1(n71), .A2(n3), .ZN(\U3/U1/Z_3 ) );
  CKND2D0 U91 ( .A1(mantissa_shift[3]), .A2(n72), .ZN(n3) );
  NR2D0 U92 ( .A1(n71), .A2(n1), .ZN(\U3/U1/Z_2 ) );
  CKND2D0 U93 ( .A1(mantissa_shift[2]), .A2(n72), .ZN(n1) );
  NR2D0 U94 ( .A1(n71), .A2(n2), .ZN(\U3/U1/Z_1 ) );
  CKND2D0 U95 ( .A1(mantissa_shift[1]), .A2(n72), .ZN(n2) );
  CKND0 U96 ( .I(\U3/U2/Z_0 ), .ZN(n71) );
  AO21D0 U97 ( .A1(\U3/U2/Z_0 ), .A2(N11), .B(mantissa_ab_c_in[21]), .Z(
        \U3/U1/Z_0 ) );
  NR2D0 U98 ( .A1(mantissa_ab_c_in[20]), .A2(mantissa_ab_c_in[21]), .ZN(
        \U3/U2/Z_0 ) );
  AN2D0 U99 ( .A1(mantissa_shift[0]), .A2(n72), .Z(N11) );
  AN4D0 U100 ( .A1(exp_ab_c_in[4]), .A2(exp_ab_c_in[3]), .A3(n73), .A4(
        exp_ab_c_in[2]), .Z(n72) );
  AN2D0 U101 ( .A1(exp_ab_c_in[0]), .A2(exp_ab_c_in[1]), .Z(n73) );
endmodule


module fma_top_1 ( a, b, c, fma_en, clk, rst, z, fma_vld );
  input [15:0] a;
  input [15:0] b;
  input [15:0] c;
  output [15:0] z;
  input fma_en, clk, rst;
  output fma_vld;
  wire   N4, a_equals_one, b_equals_one, fma_en_ff, exp_ab_greater,
         exp_ab_less, exp_diff_done, sign_ab, mult_done, adder_done, _0_net_,
         rounder_done, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;
  wire   [15:0] a_ff;
  wire   [15:0] b_ff;
  wire   [15:0] c_ff;
  wire   [4:0] exp_diff;
  wire   [4:0] exp_ab;
  wire   [19:0] mantissa_ab;
  wire   [21:0] mantissa_ab_c;
  wire   [4:0] exp_ab_c;
  wire   [15:0] result;
  wire   [4:0] mantissa_shift;
  wire   [4:0] exp_ab_c_out;
  tri   rst;
  assign fma_vld = rounder_done;

  fma_exp_diff_1 fma_exp_diff_i ( .exp_a(a_ff[14:10]), .exp_b(b_ff[14:10]), 
        .exp_c(c_ff[14:10]), .exp_diff_start(fma_en_ff), .fma_byp(N4), 
        .exp_diff(exp_diff), .exp_ab(exp_ab), .exp_ab_greater(exp_ab_greater), 
        .exp_ab_less(exp_ab_less), .exp_diff_done(exp_diff_done) );
  fma_mult_tree_1 fma_mult_tree_i ( .mantissa_a(a_ff[9:0]), .mantissa_b(
        b_ff[9:0]), .sign_a(a_ff[15]), .sign_b(b_ff[15]), .fma_byp(N4), 
        .a_equals_one(a_equals_one), .b_equals_one(b_equals_one), .mult_start(
        fma_en_ff), .mantissa_ab(mantissa_ab), .sign_ab(sign_ab), .mult_done(
        mult_done) );
  fma_aligner_adder_1 fma_aligner_adder_i ( .mantissa_ab(mantissa_ab), 
        .exp_ab(exp_ab), .sign_ab(sign_ab), .c(c_ff), .exp_diff(exp_diff), 
        .exp_ab_greater(exp_ab_greater), .exp_ab_less(exp_ab_less), .fma_byp(
        N4), .add_byp(n31), .adder_start(_0_net_), .mantissa_ab_c(
        mantissa_ab_c), .exp_ab_c(exp_ab_c), .sign_ab_c(result[15]), 
        .mantissa_shift(mantissa_shift), .adder_done(adder_done) );
  fma_normalizer_rounder_1 fma_normalizer_rounder_i ( .mantissa_ab_c_in(
        mantissa_ab_c), .exp_ab_c_in(exp_ab_c), .mantissa_shift(mantissa_shift), .fma_byp(N4), .rounder_start(adder_done), .mantissa_ab_c_out(result[9:0]), 
        .exp_ab_c_out(exp_ab_c_out), .rounder_done(rounder_done) );
  DFKCNQD1 \a_ff_reg[15]  ( .CN(n30), .D(a[15]), .CP(clk), .Q(a_ff[15]) );
  DFKCNQD1 \b_ff_reg[10]  ( .CN(n30), .D(b[10]), .CP(clk), .Q(b_ff[10]) );
  DFKCNQD1 \a_ff_reg[14]  ( .CN(n30), .D(a[14]), .CP(clk), .Q(a_ff[14]) );
  DFKCNQD1 \a_ff_reg[10]  ( .CN(n30), .D(a[10]), .CP(clk), .Q(a_ff[10]) );
  DFKCNQD1 \b_ff_reg[14]  ( .CN(n30), .D(b[14]), .CP(clk), .Q(b_ff[14]) );
  DFKCNQD1 \b_ff_reg[8]  ( .CN(n30), .D(b[8]), .CP(clk), .Q(b_ff[8]) );
  DFKCNQD1 \b_ff_reg[15]  ( .CN(n30), .D(b[15]), .CP(clk), .Q(b_ff[15]) );
  DFKCNQD1 \b_ff_reg[11]  ( .CN(n30), .D(b[11]), .CP(clk), .Q(b_ff[11]) );
  DFKCNQD1 \a_ff_reg[12]  ( .CN(n30), .D(a[12]), .CP(clk), .Q(a_ff[12]) );
  DFKCNQD1 \b_ff_reg[12]  ( .CN(n30), .D(b[12]), .CP(clk), .Q(b_ff[12]) );
  DFKCNQD1 \c_ff_reg[5]  ( .CN(n30), .D(c[5]), .CP(clk), .Q(c_ff[5]) );
  DFKCNQD1 \a_ff_reg[13]  ( .CN(n30), .D(a[13]), .CP(clk), .Q(a_ff[13]) );
  DFKCNQD1 \a_ff_reg[11]  ( .CN(n30), .D(a[11]), .CP(clk), .Q(a_ff[11]) );
  DFKCNQD1 \b_ff_reg[13]  ( .CN(n30), .D(b[13]), .CP(clk), .Q(b_ff[13]) );
  DFKCNQD1 \c_ff_reg[8]  ( .CN(n30), .D(c[8]), .CP(clk), .Q(c_ff[8]) );
  DFKCNQD1 \b_ff_reg[4]  ( .CN(n30), .D(b[4]), .CP(clk), .Q(b_ff[4]) );
  DFKCNQD1 \b_ff_reg[2]  ( .CN(n30), .D(b[2]), .CP(clk), .Q(b_ff[2]) );
  DFKCNQD1 \c_ff_reg[4]  ( .CN(n30), .D(c[4]), .CP(clk), .Q(c_ff[4]) );
  DFKCNQD1 \b_ff_reg[6]  ( .CN(n30), .D(b[6]), .CP(clk), .Q(b_ff[6]) );
  DFKCNQD1 \c_ff_reg[10]  ( .CN(n30), .D(c[10]), .CP(clk), .Q(c_ff[10]) );
  DFKCNQD1 \c_ff_reg[9]  ( .CN(n30), .D(c[9]), .CP(clk), .Q(c_ff[9]) );
  DFKCNQD1 \c_ff_reg[12]  ( .CN(n30), .D(c[12]), .CP(clk), .Q(c_ff[12]) );
  DFKCNQD1 \c_ff_reg[14]  ( .CN(n30), .D(c[14]), .CP(clk), .Q(c_ff[14]) );
  DFKCNQD1 \c_ff_reg[13]  ( .CN(n30), .D(c[13]), .CP(clk), .Q(c_ff[13]) );
  DFKCNQD1 \c_ff_reg[3]  ( .CN(n30), .D(c[3]), .CP(clk), .Q(c_ff[3]) );
  DFKCNQD1 \c_ff_reg[1]  ( .CN(n30), .D(c[1]), .CP(clk), .Q(c_ff[1]) );
  DFKCNQD1 \c_ff_reg[7]  ( .CN(n30), .D(c[7]), .CP(clk), .Q(c_ff[7]) );
  DFKCNQD1 \c_ff_reg[0]  ( .CN(n30), .D(c[0]), .CP(clk), .Q(c_ff[0]) );
  DFKCNQD1 \b_ff_reg[1]  ( .CN(n30), .D(b[1]), .CP(clk), .Q(b_ff[1]) );
  DFKCNQD1 \c_ff_reg[2]  ( .CN(n30), .D(c[2]), .CP(clk), .Q(c_ff[2]) );
  DFKCNQD1 \c_ff_reg[6]  ( .CN(n30), .D(c[6]), .CP(clk), .Q(c_ff[6]) );
  DFKCNQD1 \c_ff_reg[11]  ( .CN(n30), .D(c[11]), .CP(clk), .Q(c_ff[11]) );
  DFKCNQD1 \a_ff_reg[9]  ( .CN(n30), .D(a[9]), .CP(clk), .Q(a_ff[9]) );
  DFKCNQD1 \b_ff_reg[3]  ( .CN(n30), .D(b[3]), .CP(clk), .Q(b_ff[3]) );
  DFKCNQD1 \a_ff_reg[0]  ( .CN(n30), .D(a[0]), .CP(clk), .Q(a_ff[0]) );
  DFKCNQD1 \c_ff_reg[15]  ( .CN(n30), .D(c[15]), .CP(clk), .Q(c_ff[15]) );
  DFKCNQD1 \b_ff_reg[5]  ( .CN(n30), .D(b[5]), .CP(clk), .Q(b_ff[5]) );
  DFKCNQD1 \a_ff_reg[7]  ( .CN(n30), .D(a[7]), .CP(clk), .Q(a_ff[7]) );
  DFKCNQD1 \b_ff_reg[0]  ( .CN(n30), .D(b[0]), .CP(clk), .Q(b_ff[0]) );
  DFKCNQD1 \a_ff_reg[4]  ( .CN(n30), .D(a[4]), .CP(clk), .Q(a_ff[4]) );
  DFKCNQD1 \a_ff_reg[8]  ( .CN(n30), .D(a[8]), .CP(clk), .Q(a_ff[8]) );
  DFKCNQD1 \a_ff_reg[1]  ( .CN(n30), .D(a[1]), .CP(clk), .Q(a_ff[1]) );
  DFKCNQD1 \a_ff_reg[3]  ( .CN(n30), .D(a[3]), .CP(clk), .Q(a_ff[3]) );
  DFKCNQD1 \a_ff_reg[5]  ( .CN(n30), .D(a[5]), .CP(clk), .Q(a_ff[5]) );
  DFKCNQD1 \a_ff_reg[2]  ( .CN(n30), .D(a[2]), .CP(clk), .Q(a_ff[2]) );
  DFKCNQD1 \a_ff_reg[6]  ( .CN(n30), .D(a[6]), .CP(clk), .Q(a_ff[6]) );
  DFKCNQD1 \b_ff_reg[7]  ( .CN(n30), .D(b[7]), .CP(clk), .Q(b_ff[7]) );
  DFKCNQD1 \b_ff_reg[9]  ( .CN(n30), .D(b[9]), .CP(clk), .Q(b_ff[9]) );
  DFKCNQD1 fma_en_ff_reg ( .CN(n30), .D(fma_en), .CP(clk), .Q(fma_en_ff) );
  INVD1 U3 ( .I(rst), .ZN(n30) );
  ND2D1 U4 ( .A1(n18), .A2(n19), .ZN(N4) );
  TIEL U5 ( .ZN(z[15]) );
  AN2D0 U6 ( .A1(result[9]), .A2(n1), .Z(z[9]) );
  AN2D0 U7 ( .A1(result[8]), .A2(n1), .Z(z[8]) );
  AN2D0 U8 ( .A1(result[7]), .A2(n1), .Z(z[7]) );
  AN2D0 U9 ( .A1(result[6]), .A2(n1), .Z(z[6]) );
  AN2D0 U10 ( .A1(result[5]), .A2(n1), .Z(z[5]) );
  AN2D0 U11 ( .A1(result[4]), .A2(n1), .Z(z[4]) );
  AN2D0 U12 ( .A1(result[3]), .A2(n1), .Z(z[3]) );
  AN2D0 U13 ( .A1(result[2]), .A2(n1), .Z(z[2]) );
  AN2D0 U14 ( .A1(result[1]), .A2(n1), .Z(z[1]) );
  IOA21D0 U15 ( .A1(exp_ab_c_out[4]), .A2(n1), .B(n2), .ZN(z[14]) );
  IOA21D0 U16 ( .A1(exp_ab_c_out[3]), .A2(n1), .B(n2), .ZN(z[13]) );
  IOA21D0 U17 ( .A1(exp_ab_c_out[2]), .A2(n1), .B(n2), .ZN(z[12]) );
  IOA21D0 U18 ( .A1(exp_ab_c_out[1]), .A2(n1), .B(n2), .ZN(z[11]) );
  IOA21D0 U19 ( .A1(exp_ab_c_out[0]), .A2(n1), .B(n2), .ZN(z[10]) );
  OR2D0 U20 ( .A1(n3), .A2(result[15]), .Z(n2) );
  AOI33D0 U21 ( .A1(c_ff[14]), .A2(c_ff[13]), .A3(n4), .B1(exp_ab[4]), .B2(
        exp_ab[3]), .B3(n5), .ZN(n3) );
  AN3D0 U22 ( .A1(exp_ab[1]), .A2(exp_ab[0]), .A3(exp_ab[2]), .Z(n5) );
  AN3D0 U23 ( .A1(c_ff[12]), .A2(c_ff[10]), .A3(c_ff[11]), .Z(n4) );
  AN2D0 U24 ( .A1(result[0]), .A2(n1), .Z(z[0]) );
  CKND0 U25 ( .I(result[15]), .ZN(n1) );
  AN4D0 U26 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n31) );
  NR4D0 U27 ( .A1(c_ff[9]), .A2(c_ff[8]), .A3(c_ff[7]), .A4(c_ff[6]), .ZN(n9)
         );
  NR4D0 U28 ( .A1(c_ff[5]), .A2(c_ff[4]), .A3(c_ff[3]), .A4(c_ff[2]), .ZN(n8)
         );
  NR4D0 U29 ( .A1(c_ff[1]), .A2(c_ff[14]), .A3(c_ff[13]), .A4(c_ff[12]), .ZN(
        n7) );
  NR3D0 U30 ( .A1(c_ff[0]), .A2(c_ff[11]), .A3(c_ff[10]), .ZN(n6) );
  NR4D0 U31 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(b_equals_one) );
  CKND2D0 U32 ( .A1(b_ff[13]), .A2(b_ff[12]), .ZN(n10) );
  NR4D0 U33 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(a_equals_one) );
  CKND2D0 U34 ( .A1(a_ff[13]), .A2(a_ff[12]), .ZN(n14) );
  AN2D0 U35 ( .A1(mult_done), .A2(exp_diff_done), .Z(_0_net_) );
  IND4D0 U36 ( .A1(n16), .B1(n17), .B2(n15), .B3(n20), .ZN(n19) );
  NR3D0 U37 ( .A1(a_ff[12]), .A2(a_ff[15]), .A3(a_ff[13]), .ZN(n20) );
  CKND0 U38 ( .I(a_ff[11]), .ZN(n15) );
  CKND0 U39 ( .I(a_ff[10]), .ZN(n17) );
  ND4D0 U40 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n16) );
  NR3D0 U41 ( .A1(a_ff[7]), .A2(a_ff[9]), .A3(a_ff[8]), .ZN(n24) );
  NR3D0 U42 ( .A1(a_ff[4]), .A2(a_ff[6]), .A3(a_ff[5]), .ZN(n23) );
  NR3D0 U43 ( .A1(a_ff[1]), .A2(a_ff[3]), .A3(a_ff[2]), .ZN(n22) );
  NR2D0 U44 ( .A1(a_ff[14]), .A2(a_ff[0]), .ZN(n21) );
  IND4D0 U45 ( .A1(n12), .B1(n13), .B2(n11), .B3(n25), .ZN(n18) );
  NR3D0 U46 ( .A1(b_ff[12]), .A2(b_ff[15]), .A3(b_ff[13]), .ZN(n25) );
  CKND0 U47 ( .I(b_ff[11]), .ZN(n11) );
  CKND0 U48 ( .I(b_ff[10]), .ZN(n13) );
  ND4D0 U49 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n12) );
  NR3D0 U50 ( .A1(b_ff[7]), .A2(b_ff[9]), .A3(b_ff[8]), .ZN(n29) );
  NR3D0 U51 ( .A1(b_ff[4]), .A2(b_ff[6]), .A3(b_ff[5]), .ZN(n28) );
  NR3D0 U52 ( .A1(b_ff[1]), .A2(b_ff[3]), .A3(b_ff[2]), .ZN(n27) );
  NR2D0 U53 ( .A1(b_ff[14]), .A2(b_ff[0]), .ZN(n26) );
endmodule


module neuron_1 ( input_value, input_weight, input_bias, rst, en, srdy, 
        output_value, drdy, done, clk );
  input [127:0] input_value;
  input [127:0] input_weight;
  input [15:0] input_bias;
  output [15:0] output_value;
  input rst, en, srdy, clk;
  output drdy, done;
  wire   \*Logic1* , \input_value_loc[7][15] , \input_value_loc[7][14] ,
         \input_value_loc[7][13] , \input_value_loc[7][12] ,
         \input_value_loc[7][11] , \input_value_loc[7][10] ,
         \input_value_loc[7][9] , \input_value_loc[7][8] ,
         \input_value_loc[7][7] , \input_value_loc[7][6] ,
         \input_value_loc[7][5] , \input_value_loc[7][4] ,
         \input_value_loc[7][3] , \input_value_loc[7][2] ,
         \input_value_loc[7][1] , \input_value_loc[7][0] ,
         \input_value_loc[6][15] , \input_value_loc[6][14] ,
         \input_value_loc[6][13] , \input_value_loc[6][12] ,
         \input_value_loc[6][11] , \input_value_loc[6][10] ,
         \input_value_loc[6][9] , \input_value_loc[6][8] ,
         \input_value_loc[6][7] , \input_value_loc[6][6] ,
         \input_value_loc[6][5] , \input_value_loc[6][4] ,
         \input_value_loc[6][3] , \input_value_loc[6][2] ,
         \input_value_loc[6][1] , \input_value_loc[6][0] ,
         \input_value_loc[5][15] , \input_value_loc[5][14] ,
         \input_value_loc[5][13] , \input_value_loc[5][12] ,
         \input_value_loc[5][11] , \input_value_loc[5][10] ,
         \input_value_loc[5][9] , \input_value_loc[5][8] ,
         \input_value_loc[5][7] , \input_value_loc[5][6] ,
         \input_value_loc[5][5] , \input_value_loc[5][4] ,
         \input_value_loc[5][3] , \input_value_loc[5][2] ,
         \input_value_loc[5][1] , \input_value_loc[5][0] ,
         \input_value_loc[4][15] , \input_value_loc[4][14] ,
         \input_value_loc[4][13] , \input_value_loc[4][12] ,
         \input_value_loc[4][11] , \input_value_loc[4][10] ,
         \input_value_loc[4][9] , \input_value_loc[4][8] ,
         \input_value_loc[4][7] , \input_value_loc[4][6] ,
         \input_value_loc[4][5] , \input_value_loc[4][4] ,
         \input_value_loc[4][3] , \input_value_loc[4][2] ,
         \input_value_loc[4][1] , \input_value_loc[4][0] ,
         \input_value_loc[3][15] , \input_value_loc[3][14] ,
         \input_value_loc[3][13] , \input_value_loc[3][12] ,
         \input_value_loc[3][11] , \input_value_loc[3][10] ,
         \input_value_loc[3][9] , \input_value_loc[3][8] ,
         \input_value_loc[3][7] , \input_value_loc[3][6] ,
         \input_value_loc[3][5] , \input_value_loc[3][4] ,
         \input_value_loc[3][3] , \input_value_loc[3][2] ,
         \input_value_loc[3][1] , \input_value_loc[3][0] ,
         \input_value_loc[2][15] , \input_value_loc[2][14] ,
         \input_value_loc[2][13] , \input_value_loc[2][12] ,
         \input_value_loc[2][11] , \input_value_loc[2][10] ,
         \input_value_loc[2][9] , \input_value_loc[2][8] ,
         \input_value_loc[2][7] , \input_value_loc[2][6] ,
         \input_value_loc[2][5] , \input_value_loc[2][4] ,
         \input_value_loc[2][3] , \input_value_loc[2][2] ,
         \input_value_loc[2][1] , \input_value_loc[2][0] ,
         \input_value_loc[1][15] , \input_value_loc[1][14] ,
         \input_value_loc[1][13] , \input_value_loc[1][12] ,
         \input_value_loc[1][11] , \input_value_loc[1][10] ,
         \input_value_loc[1][9] , \input_value_loc[1][8] ,
         \input_value_loc[1][7] , \input_value_loc[1][6] ,
         \input_value_loc[1][5] , \input_value_loc[1][4] ,
         \input_value_loc[1][3] , \input_value_loc[1][2] ,
         \input_value_loc[1][1] , \input_value_loc[1][0] ,
         \input_value_loc[0][15] , \input_value_loc[0][14] ,
         \input_value_loc[0][13] , \input_value_loc[0][12] ,
         \input_value_loc[0][11] , \input_value_loc[0][10] ,
         \input_value_loc[0][9] , \input_value_loc[0][8] ,
         \input_value_loc[0][7] , \input_value_loc[0][6] ,
         \input_value_loc[0][5] , \input_value_loc[0][4] ,
         \input_value_loc[0][3] , \input_value_loc[0][2] ,
         \input_value_loc[0][1] , \input_value_loc[0][0] ,
         \input_weight_loc[7][15] , \input_weight_loc[7][14] ,
         \input_weight_loc[7][13] , \input_weight_loc[7][12] ,
         \input_weight_loc[7][11] , \input_weight_loc[7][10] ,
         \input_weight_loc[7][9] , \input_weight_loc[7][8] ,
         \input_weight_loc[7][7] , \input_weight_loc[7][6] ,
         \input_weight_loc[7][5] , \input_weight_loc[7][4] ,
         \input_weight_loc[7][3] , \input_weight_loc[7][2] ,
         \input_weight_loc[7][1] , \input_weight_loc[7][0] ,
         \input_weight_loc[6][15] , \input_weight_loc[6][14] ,
         \input_weight_loc[6][13] , \input_weight_loc[6][12] ,
         \input_weight_loc[6][11] , \input_weight_loc[6][10] ,
         \input_weight_loc[6][9] , \input_weight_loc[6][8] ,
         \input_weight_loc[6][7] , \input_weight_loc[6][6] ,
         \input_weight_loc[6][5] , \input_weight_loc[6][4] ,
         \input_weight_loc[6][3] , \input_weight_loc[6][2] ,
         \input_weight_loc[6][1] , \input_weight_loc[6][0] ,
         \input_weight_loc[5][15] , \input_weight_loc[5][14] ,
         \input_weight_loc[5][13] , \input_weight_loc[5][12] ,
         \input_weight_loc[5][11] , \input_weight_loc[5][10] ,
         \input_weight_loc[5][9] , \input_weight_loc[5][8] ,
         \input_weight_loc[5][7] , \input_weight_loc[5][6] ,
         \input_weight_loc[5][5] , \input_weight_loc[5][4] ,
         \input_weight_loc[5][3] , \input_weight_loc[5][2] ,
         \input_weight_loc[5][1] , \input_weight_loc[5][0] ,
         \input_weight_loc[4][15] , \input_weight_loc[4][14] ,
         \input_weight_loc[4][13] , \input_weight_loc[4][12] ,
         \input_weight_loc[4][11] , \input_weight_loc[4][10] ,
         \input_weight_loc[4][9] , \input_weight_loc[4][8] ,
         \input_weight_loc[4][7] , \input_weight_loc[4][6] ,
         \input_weight_loc[4][5] , \input_weight_loc[4][4] ,
         \input_weight_loc[4][3] , \input_weight_loc[4][2] ,
         \input_weight_loc[4][1] , \input_weight_loc[4][0] ,
         \input_weight_loc[3][15] , \input_weight_loc[3][14] ,
         \input_weight_loc[3][13] , \input_weight_loc[3][12] ,
         \input_weight_loc[3][11] , \input_weight_loc[3][10] ,
         \input_weight_loc[3][9] , \input_weight_loc[3][8] ,
         \input_weight_loc[3][7] , \input_weight_loc[3][6] ,
         \input_weight_loc[3][5] , \input_weight_loc[3][4] ,
         \input_weight_loc[3][3] , \input_weight_loc[3][2] ,
         \input_weight_loc[3][1] , \input_weight_loc[3][0] ,
         \input_weight_loc[2][15] , \input_weight_loc[2][14] ,
         \input_weight_loc[2][13] , \input_weight_loc[2][12] ,
         \input_weight_loc[2][11] , \input_weight_loc[2][10] ,
         \input_weight_loc[2][9] , \input_weight_loc[2][8] ,
         \input_weight_loc[2][7] , \input_weight_loc[2][6] ,
         \input_weight_loc[2][5] , \input_weight_loc[2][4] ,
         \input_weight_loc[2][3] , \input_weight_loc[2][2] ,
         \input_weight_loc[2][1] , \input_weight_loc[2][0] ,
         \input_weight_loc[1][15] , \input_weight_loc[1][14] ,
         \input_weight_loc[1][13] , \input_weight_loc[1][12] ,
         \input_weight_loc[1][11] , \input_weight_loc[1][10] ,
         \input_weight_loc[1][9] , \input_weight_loc[1][8] ,
         \input_weight_loc[1][7] , \input_weight_loc[1][6] ,
         \input_weight_loc[1][5] , \input_weight_loc[1][4] ,
         \input_weight_loc[1][3] , \input_weight_loc[1][2] ,
         \input_weight_loc[1][1] , \input_weight_loc[1][0] ,
         \input_weight_loc[0][15] , \input_weight_loc[0][14] ,
         \input_weight_loc[0][13] , \input_weight_loc[0][12] ,
         \input_weight_loc[0][11] , \input_weight_loc[0][10] ,
         \input_weight_loc[0][9] , \input_weight_loc[0][8] ,
         \input_weight_loc[0][7] , \input_weight_loc[0][6] ,
         \input_weight_loc[0][5] , \input_weight_loc[0][4] ,
         \input_weight_loc[0][3] , \input_weight_loc[0][2] ,
         \input_weight_loc[0][1] , \input_weight_loc[0][0] , N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150;
  wire   [3:0] cur_state;
  wire   [3:0] nxt_state;
  wire   [15:0] fma_a;
  wire   [15:0] fma_b;
  wire   [15:0] output_value_loc;
  wire   [15:0] fma_z;
  tri   rst;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign done = \*Logic1* ;
  assign drdy = \*Logic1* ;

  LHQD1 \fma_a_reg[0]  ( .E(N90), .D(N91), .Q(fma_a[0]) );
  LHQD1 \fma_a_reg[1]  ( .E(N90), .D(N92), .Q(fma_a[1]) );
  LHQD1 \fma_a_reg[2]  ( .E(N90), .D(N93), .Q(fma_a[2]) );
  LHQD1 \fma_a_reg[3]  ( .E(N90), .D(N94), .Q(fma_a[3]) );
  LHQD1 \fma_a_reg[4]  ( .E(N90), .D(N95), .Q(fma_a[4]) );
  LHQD1 \fma_a_reg[5]  ( .E(N90), .D(N96), .Q(fma_a[5]) );
  LHQD1 \fma_a_reg[6]  ( .E(N90), .D(N97), .Q(fma_a[6]) );
  LHQD1 \fma_a_reg[7]  ( .E(N90), .D(N98), .Q(fma_a[7]) );
  LHQD1 \fma_a_reg[8]  ( .E(N90), .D(N99), .Q(fma_a[8]) );
  LHQD1 \fma_a_reg[15]  ( .E(N90), .D(N106), .Q(fma_a[15]) );
  LHQD1 \fma_a_reg[14]  ( .E(N90), .D(N105), .Q(fma_a[14]) );
  LHQD1 \fma_a_reg[13]  ( .E(N90), .D(N104), .Q(fma_a[13]) );
  LHQD1 \fma_a_reg[12]  ( .E(N90), .D(N103), .Q(fma_a[12]) );
  LHQD1 \fma_a_reg[11]  ( .E(N90), .D(N102), .Q(fma_a[11]) );
  LHQD1 \fma_a_reg[10]  ( .E(N90), .D(N101), .Q(fma_a[10]) );
  LHQD1 \fma_a_reg[9]  ( .E(N90), .D(N100), .Q(fma_a[9]) );
  LHQD1 \fma_b_reg[0]  ( .E(N90), .D(N107), .Q(fma_b[0]) );
  LHQD1 \fma_b_reg[1]  ( .E(N90), .D(N108), .Q(fma_b[1]) );
  LHQD1 \fma_b_reg[2]  ( .E(N90), .D(N109), .Q(fma_b[2]) );
  LHQD1 \fma_b_reg[3]  ( .E(N90), .D(N110), .Q(fma_b[3]) );
  LHQD1 \fma_b_reg[4]  ( .E(N90), .D(N111), .Q(fma_b[4]) );
  LHQD1 \fma_b_reg[5]  ( .E(N90), .D(N112), .Q(fma_b[5]) );
  LHQD1 \fma_b_reg[6]  ( .E(N90), .D(N113), .Q(fma_b[6]) );
  LHQD1 \fma_b_reg[7]  ( .E(N90), .D(N114), .Q(fma_b[7]) );
  LHQD1 \fma_b_reg[8]  ( .E(N90), .D(N115), .Q(fma_b[8]) );
  LHQD1 \fma_b_reg[9]  ( .E(N90), .D(N116), .Q(fma_b[9]) );
  LHQD1 \fma_b_reg[10]  ( .E(N90), .D(N117), .Q(fma_b[10]) );
  LHQD1 \fma_b_reg[11]  ( .E(N90), .D(N118), .Q(fma_b[11]) );
  LHQD1 \fma_b_reg[12]  ( .E(N90), .D(N119), .Q(fma_b[12]) );
  LHQD1 \fma_b_reg[13]  ( .E(N90), .D(N120), .Q(fma_b[13]) );
  LHQD1 \fma_b_reg[14]  ( .E(N90), .D(N121), .Q(fma_b[14]) );
  LHQD1 \fma_b_reg[15]  ( .E(N90), .D(N122), .Q(fma_b[15]) );
  fma_top_1 u_neuron ( .a(fma_a), .b(fma_b), .c({n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1}), .fma_en(\*Logic1* ), .clk(clk), 
        .rst(rst), .z({SYNOPSYS_UNCONNECTED__0, fma_z[14:0]}) );
  DFQD1 \input_weight_loc_reg[6][15]  ( .D(input_weight[31]), .CP(srdy), .Q(
        \input_weight_loc[6][15] ) );
  DFQD1 \input_weight_loc_reg[6][14]  ( .D(input_weight[30]), .CP(srdy), .Q(
        \input_weight_loc[6][14] ) );
  DFQD1 \input_weight_loc_reg[6][13]  ( .D(input_weight[29]), .CP(srdy), .Q(
        \input_weight_loc[6][13] ) );
  DFQD1 \input_weight_loc_reg[6][12]  ( .D(input_weight[28]), .CP(srdy), .Q(
        \input_weight_loc[6][12] ) );
  DFQD1 \input_weight_loc_reg[6][11]  ( .D(input_weight[27]), .CP(srdy), .Q(
        \input_weight_loc[6][11] ) );
  DFQD1 \input_weight_loc_reg[6][10]  ( .D(input_weight[26]), .CP(srdy), .Q(
        \input_weight_loc[6][10] ) );
  DFQD1 \input_weight_loc_reg[6][9]  ( .D(input_weight[25]), .CP(srdy), .Q(
        \input_weight_loc[6][9] ) );
  DFQD1 \input_weight_loc_reg[6][8]  ( .D(input_weight[24]), .CP(srdy), .Q(
        \input_weight_loc[6][8] ) );
  DFQD1 \input_weight_loc_reg[6][7]  ( .D(input_weight[23]), .CP(srdy), .Q(
        \input_weight_loc[6][7] ) );
  DFQD1 \input_weight_loc_reg[6][6]  ( .D(input_weight[22]), .CP(srdy), .Q(
        \input_weight_loc[6][6] ) );
  DFQD1 \input_weight_loc_reg[6][5]  ( .D(input_weight[21]), .CP(srdy), .Q(
        \input_weight_loc[6][5] ) );
  DFQD1 \input_weight_loc_reg[6][4]  ( .D(input_weight[20]), .CP(srdy), .Q(
        \input_weight_loc[6][4] ) );
  DFQD1 \input_weight_loc_reg[6][3]  ( .D(input_weight[19]), .CP(srdy), .Q(
        \input_weight_loc[6][3] ) );
  DFQD1 \input_weight_loc_reg[6][2]  ( .D(input_weight[18]), .CP(srdy), .Q(
        \input_weight_loc[6][2] ) );
  DFQD1 \input_weight_loc_reg[6][1]  ( .D(input_weight[17]), .CP(srdy), .Q(
        \input_weight_loc[6][1] ) );
  DFQD1 \input_weight_loc_reg[6][0]  ( .D(input_weight[16]), .CP(srdy), .Q(
        \input_weight_loc[6][0] ) );
  DFQD1 \input_weight_loc_reg[3][15]  ( .D(input_weight[79]), .CP(srdy), .Q(
        \input_weight_loc[3][15] ) );
  DFQD1 \input_weight_loc_reg[3][14]  ( .D(input_weight[78]), .CP(srdy), .Q(
        \input_weight_loc[3][14] ) );
  DFQD1 \input_weight_loc_reg[3][13]  ( .D(input_weight[77]), .CP(srdy), .Q(
        \input_weight_loc[3][13] ) );
  DFQD1 \input_weight_loc_reg[3][12]  ( .D(input_weight[76]), .CP(srdy), .Q(
        \input_weight_loc[3][12] ) );
  DFQD1 \input_weight_loc_reg[3][11]  ( .D(input_weight[75]), .CP(srdy), .Q(
        \input_weight_loc[3][11] ) );
  DFQD1 \input_weight_loc_reg[3][10]  ( .D(input_weight[74]), .CP(srdy), .Q(
        \input_weight_loc[3][10] ) );
  DFQD1 \input_weight_loc_reg[3][9]  ( .D(input_weight[73]), .CP(srdy), .Q(
        \input_weight_loc[3][9] ) );
  DFQD1 \input_weight_loc_reg[3][8]  ( .D(input_weight[72]), .CP(srdy), .Q(
        \input_weight_loc[3][8] ) );
  DFQD1 \input_weight_loc_reg[3][7]  ( .D(input_weight[71]), .CP(srdy), .Q(
        \input_weight_loc[3][7] ) );
  DFQD1 \input_weight_loc_reg[3][6]  ( .D(input_weight[70]), .CP(srdy), .Q(
        \input_weight_loc[3][6] ) );
  DFQD1 \input_weight_loc_reg[3][5]  ( .D(input_weight[69]), .CP(srdy), .Q(
        \input_weight_loc[3][5] ) );
  DFQD1 \input_weight_loc_reg[3][4]  ( .D(input_weight[68]), .CP(srdy), .Q(
        \input_weight_loc[3][4] ) );
  DFQD1 \input_weight_loc_reg[3][3]  ( .D(input_weight[67]), .CP(srdy), .Q(
        \input_weight_loc[3][3] ) );
  DFQD1 \input_weight_loc_reg[3][2]  ( .D(input_weight[66]), .CP(srdy), .Q(
        \input_weight_loc[3][2] ) );
  DFQD1 \input_weight_loc_reg[3][1]  ( .D(input_weight[65]), .CP(srdy), .Q(
        \input_weight_loc[3][1] ) );
  DFQD1 \input_weight_loc_reg[3][0]  ( .D(input_weight[64]), .CP(srdy), .Q(
        \input_weight_loc[3][0] ) );
  DFQD1 \input_weight_loc_reg[1][15]  ( .D(input_weight[111]), .CP(srdy), .Q(
        \input_weight_loc[1][15] ) );
  DFQD1 \input_weight_loc_reg[1][14]  ( .D(input_weight[110]), .CP(srdy), .Q(
        \input_weight_loc[1][14] ) );
  DFQD1 \input_weight_loc_reg[1][13]  ( .D(input_weight[109]), .CP(srdy), .Q(
        \input_weight_loc[1][13] ) );
  DFQD1 \input_weight_loc_reg[1][12]  ( .D(input_weight[108]), .CP(srdy), .Q(
        \input_weight_loc[1][12] ) );
  DFQD1 \input_weight_loc_reg[1][11]  ( .D(input_weight[107]), .CP(srdy), .Q(
        \input_weight_loc[1][11] ) );
  DFQD1 \input_weight_loc_reg[1][10]  ( .D(input_weight[106]), .CP(srdy), .Q(
        \input_weight_loc[1][10] ) );
  DFQD1 \input_weight_loc_reg[1][9]  ( .D(input_weight[105]), .CP(srdy), .Q(
        \input_weight_loc[1][9] ) );
  DFQD1 \input_weight_loc_reg[1][8]  ( .D(input_weight[104]), .CP(srdy), .Q(
        \input_weight_loc[1][8] ) );
  DFQD1 \input_weight_loc_reg[1][7]  ( .D(input_weight[103]), .CP(srdy), .Q(
        \input_weight_loc[1][7] ) );
  DFQD1 \input_weight_loc_reg[1][6]  ( .D(input_weight[102]), .CP(srdy), .Q(
        \input_weight_loc[1][6] ) );
  DFQD1 \input_weight_loc_reg[1][5]  ( .D(input_weight[101]), .CP(srdy), .Q(
        \input_weight_loc[1][5] ) );
  DFQD1 \input_weight_loc_reg[1][4]  ( .D(input_weight[100]), .CP(srdy), .Q(
        \input_weight_loc[1][4] ) );
  DFQD1 \input_weight_loc_reg[1][3]  ( .D(input_weight[99]), .CP(srdy), .Q(
        \input_weight_loc[1][3] ) );
  DFQD1 \input_weight_loc_reg[1][2]  ( .D(input_weight[98]), .CP(srdy), .Q(
        \input_weight_loc[1][2] ) );
  DFQD1 \input_weight_loc_reg[1][1]  ( .D(input_weight[97]), .CP(srdy), .Q(
        \input_weight_loc[1][1] ) );
  DFQD1 \input_weight_loc_reg[1][0]  ( .D(input_weight[96]), .CP(srdy), .Q(
        \input_weight_loc[1][0] ) );
  DFQD1 \input_value_loc_reg[6][15]  ( .D(input_value[31]), .CP(srdy), .Q(
        \input_value_loc[6][15] ) );
  DFQD1 \input_value_loc_reg[6][14]  ( .D(input_value[30]), .CP(srdy), .Q(
        \input_value_loc[6][14] ) );
  DFQD1 \input_value_loc_reg[6][13]  ( .D(input_value[29]), .CP(srdy), .Q(
        \input_value_loc[6][13] ) );
  DFQD1 \input_value_loc_reg[6][12]  ( .D(input_value[28]), .CP(srdy), .Q(
        \input_value_loc[6][12] ) );
  DFQD1 \input_value_loc_reg[6][11]  ( .D(input_value[27]), .CP(srdy), .Q(
        \input_value_loc[6][11] ) );
  DFQD1 \input_value_loc_reg[6][10]  ( .D(input_value[26]), .CP(srdy), .Q(
        \input_value_loc[6][10] ) );
  DFQD1 \input_value_loc_reg[6][9]  ( .D(input_value[25]), .CP(srdy), .Q(
        \input_value_loc[6][9] ) );
  DFQD1 \input_value_loc_reg[6][8]  ( .D(input_value[24]), .CP(srdy), .Q(
        \input_value_loc[6][8] ) );
  DFQD1 \input_value_loc_reg[6][7]  ( .D(input_value[23]), .CP(srdy), .Q(
        \input_value_loc[6][7] ) );
  DFQD1 \input_value_loc_reg[6][6]  ( .D(input_value[22]), .CP(srdy), .Q(
        \input_value_loc[6][6] ) );
  DFQD1 \input_value_loc_reg[6][5]  ( .D(input_value[21]), .CP(srdy), .Q(
        \input_value_loc[6][5] ) );
  DFQD1 \input_value_loc_reg[6][4]  ( .D(input_value[20]), .CP(srdy), .Q(
        \input_value_loc[6][4] ) );
  DFQD1 \input_value_loc_reg[6][3]  ( .D(input_value[19]), .CP(srdy), .Q(
        \input_value_loc[6][3] ) );
  DFQD1 \input_value_loc_reg[6][2]  ( .D(input_value[18]), .CP(srdy), .Q(
        \input_value_loc[6][2] ) );
  DFQD1 \input_value_loc_reg[6][1]  ( .D(input_value[17]), .CP(srdy), .Q(
        \input_value_loc[6][1] ) );
  DFQD1 \input_value_loc_reg[6][0]  ( .D(input_value[16]), .CP(srdy), .Q(
        \input_value_loc[6][0] ) );
  DFQD1 \input_value_loc_reg[5][15]  ( .D(input_value[47]), .CP(srdy), .Q(
        \input_value_loc[5][15] ) );
  DFQD1 \input_value_loc_reg[5][14]  ( .D(input_value[46]), .CP(srdy), .Q(
        \input_value_loc[5][14] ) );
  DFQD1 \input_value_loc_reg[5][13]  ( .D(input_value[45]), .CP(srdy), .Q(
        \input_value_loc[5][13] ) );
  DFQD1 \input_value_loc_reg[5][12]  ( .D(input_value[44]), .CP(srdy), .Q(
        \input_value_loc[5][12] ) );
  DFQD1 \input_value_loc_reg[5][11]  ( .D(input_value[43]), .CP(srdy), .Q(
        \input_value_loc[5][11] ) );
  DFQD1 \input_value_loc_reg[5][10]  ( .D(input_value[42]), .CP(srdy), .Q(
        \input_value_loc[5][10] ) );
  DFQD1 \input_value_loc_reg[5][9]  ( .D(input_value[41]), .CP(srdy), .Q(
        \input_value_loc[5][9] ) );
  DFQD1 \input_value_loc_reg[5][8]  ( .D(input_value[40]), .CP(srdy), .Q(
        \input_value_loc[5][8] ) );
  DFQD1 \input_value_loc_reg[5][7]  ( .D(input_value[39]), .CP(srdy), .Q(
        \input_value_loc[5][7] ) );
  DFQD1 \input_value_loc_reg[5][6]  ( .D(input_value[38]), .CP(srdy), .Q(
        \input_value_loc[5][6] ) );
  DFQD1 \input_value_loc_reg[5][5]  ( .D(input_value[37]), .CP(srdy), .Q(
        \input_value_loc[5][5] ) );
  DFQD1 \input_value_loc_reg[5][4]  ( .D(input_value[36]), .CP(srdy), .Q(
        \input_value_loc[5][4] ) );
  DFQD1 \input_value_loc_reg[5][3]  ( .D(input_value[35]), .CP(srdy), .Q(
        \input_value_loc[5][3] ) );
  DFQD1 \input_value_loc_reg[5][2]  ( .D(input_value[34]), .CP(srdy), .Q(
        \input_value_loc[5][2] ) );
  DFQD1 \input_value_loc_reg[5][1]  ( .D(input_value[33]), .CP(srdy), .Q(
        \input_value_loc[5][1] ) );
  DFQD1 \input_value_loc_reg[3][15]  ( .D(input_value[79]), .CP(srdy), .Q(
        \input_value_loc[3][15] ) );
  DFQD1 \input_value_loc_reg[3][14]  ( .D(input_value[78]), .CP(srdy), .Q(
        \input_value_loc[3][14] ) );
  DFQD1 \input_value_loc_reg[3][13]  ( .D(input_value[77]), .CP(srdy), .Q(
        \input_value_loc[3][13] ) );
  DFQD1 \input_value_loc_reg[3][12]  ( .D(input_value[76]), .CP(srdy), .Q(
        \input_value_loc[3][12] ) );
  DFQD1 \input_value_loc_reg[3][11]  ( .D(input_value[75]), .CP(srdy), .Q(
        \input_value_loc[3][11] ) );
  DFQD1 \input_value_loc_reg[3][10]  ( .D(input_value[74]), .CP(srdy), .Q(
        \input_value_loc[3][10] ) );
  DFQD1 \input_value_loc_reg[3][9]  ( .D(input_value[73]), .CP(srdy), .Q(
        \input_value_loc[3][9] ) );
  DFQD1 \input_value_loc_reg[3][8]  ( .D(input_value[72]), .CP(srdy), .Q(
        \input_value_loc[3][8] ) );
  DFQD1 \input_value_loc_reg[3][7]  ( .D(input_value[71]), .CP(srdy), .Q(
        \input_value_loc[3][7] ) );
  DFQD1 \input_value_loc_reg[3][6]  ( .D(input_value[70]), .CP(srdy), .Q(
        \input_value_loc[3][6] ) );
  DFQD1 \input_value_loc_reg[3][5]  ( .D(input_value[69]), .CP(srdy), .Q(
        \input_value_loc[3][5] ) );
  DFQD1 \input_value_loc_reg[3][4]  ( .D(input_value[68]), .CP(srdy), .Q(
        \input_value_loc[3][4] ) );
  DFQD1 \input_value_loc_reg[3][3]  ( .D(input_value[67]), .CP(srdy), .Q(
        \input_value_loc[3][3] ) );
  DFQD1 \input_value_loc_reg[3][2]  ( .D(input_value[66]), .CP(srdy), .Q(
        \input_value_loc[3][2] ) );
  DFQD1 \input_value_loc_reg[3][1]  ( .D(input_value[65]), .CP(srdy), .Q(
        \input_value_loc[3][1] ) );
  DFQD1 \input_value_loc_reg[3][0]  ( .D(input_value[64]), .CP(srdy), .Q(
        \input_value_loc[3][0] ) );
  DFQD1 \input_value_loc_reg[1][15]  ( .D(input_value[111]), .CP(srdy), .Q(
        \input_value_loc[1][15] ) );
  DFQD1 \input_value_loc_reg[1][14]  ( .D(input_value[110]), .CP(srdy), .Q(
        \input_value_loc[1][14] ) );
  DFQD1 \input_value_loc_reg[1][13]  ( .D(input_value[109]), .CP(srdy), .Q(
        \input_value_loc[1][13] ) );
  DFQD1 \input_value_loc_reg[1][12]  ( .D(input_value[108]), .CP(srdy), .Q(
        \input_value_loc[1][12] ) );
  DFQD1 \input_value_loc_reg[1][11]  ( .D(input_value[107]), .CP(srdy), .Q(
        \input_value_loc[1][11] ) );
  DFQD1 \input_value_loc_reg[1][10]  ( .D(input_value[106]), .CP(srdy), .Q(
        \input_value_loc[1][10] ) );
  DFQD1 \input_value_loc_reg[1][9]  ( .D(input_value[105]), .CP(srdy), .Q(
        \input_value_loc[1][9] ) );
  DFQD1 \input_value_loc_reg[1][8]  ( .D(input_value[104]), .CP(srdy), .Q(
        \input_value_loc[1][8] ) );
  DFQD1 \input_value_loc_reg[1][7]  ( .D(input_value[103]), .CP(srdy), .Q(
        \input_value_loc[1][7] ) );
  DFQD1 \input_value_loc_reg[1][6]  ( .D(input_value[102]), .CP(srdy), .Q(
        \input_value_loc[1][6] ) );
  DFQD1 \input_value_loc_reg[1][5]  ( .D(input_value[101]), .CP(srdy), .Q(
        \input_value_loc[1][5] ) );
  DFQD1 \input_value_loc_reg[1][4]  ( .D(input_value[100]), .CP(srdy), .Q(
        \input_value_loc[1][4] ) );
  DFQD1 \input_value_loc_reg[1][3]  ( .D(input_value[99]), .CP(srdy), .Q(
        \input_value_loc[1][3] ) );
  DFQD1 \input_value_loc_reg[1][2]  ( .D(input_value[98]), .CP(srdy), .Q(
        \input_value_loc[1][2] ) );
  DFQD1 \input_value_loc_reg[1][1]  ( .D(input_value[97]), .CP(srdy), .Q(
        \input_value_loc[1][1] ) );
  DFQD1 \input_value_loc_reg[1][0]  ( .D(input_value[96]), .CP(srdy), .Q(
        \input_value_loc[1][0] ) );
  DFQD1 \input_weight_loc_reg[4][15]  ( .D(input_weight[63]), .CP(srdy), .Q(
        \input_weight_loc[4][15] ) );
  DFQD1 \input_weight_loc_reg[4][14]  ( .D(input_weight[62]), .CP(srdy), .Q(
        \input_weight_loc[4][14] ) );
  DFQD1 \input_weight_loc_reg[4][13]  ( .D(input_weight[61]), .CP(srdy), .Q(
        \input_weight_loc[4][13] ) );
  DFQD1 \input_weight_loc_reg[4][12]  ( .D(input_weight[60]), .CP(srdy), .Q(
        \input_weight_loc[4][12] ) );
  DFQD1 \input_weight_loc_reg[4][11]  ( .D(input_weight[59]), .CP(srdy), .Q(
        \input_weight_loc[4][11] ) );
  DFQD1 \input_weight_loc_reg[4][10]  ( .D(input_weight[58]), .CP(srdy), .Q(
        \input_weight_loc[4][10] ) );
  DFQD1 \input_weight_loc_reg[4][9]  ( .D(input_weight[57]), .CP(srdy), .Q(
        \input_weight_loc[4][9] ) );
  DFQD1 \input_weight_loc_reg[4][8]  ( .D(input_weight[56]), .CP(srdy), .Q(
        \input_weight_loc[4][8] ) );
  DFQD1 \input_weight_loc_reg[4][7]  ( .D(input_weight[55]), .CP(srdy), .Q(
        \input_weight_loc[4][7] ) );
  DFQD1 \input_weight_loc_reg[4][6]  ( .D(input_weight[54]), .CP(srdy), .Q(
        \input_weight_loc[4][6] ) );
  DFQD1 \input_weight_loc_reg[4][5]  ( .D(input_weight[53]), .CP(srdy), .Q(
        \input_weight_loc[4][5] ) );
  DFQD1 \input_weight_loc_reg[4][4]  ( .D(input_weight[52]), .CP(srdy), .Q(
        \input_weight_loc[4][4] ) );
  DFQD1 \input_weight_loc_reg[4][3]  ( .D(input_weight[51]), .CP(srdy), .Q(
        \input_weight_loc[4][3] ) );
  DFQD1 \input_weight_loc_reg[4][2]  ( .D(input_weight[50]), .CP(srdy), .Q(
        \input_weight_loc[4][2] ) );
  DFQD1 \input_weight_loc_reg[4][1]  ( .D(input_weight[49]), .CP(srdy), .Q(
        \input_weight_loc[4][1] ) );
  DFQD1 \input_weight_loc_reg[4][0]  ( .D(input_weight[48]), .CP(srdy), .Q(
        \input_weight_loc[4][0] ) );
  DFQD1 \input_weight_loc_reg[2][15]  ( .D(input_weight[95]), .CP(srdy), .Q(
        \input_weight_loc[2][15] ) );
  DFQD1 \input_weight_loc_reg[2][14]  ( .D(input_weight[94]), .CP(srdy), .Q(
        \input_weight_loc[2][14] ) );
  DFQD1 \input_weight_loc_reg[2][13]  ( .D(input_weight[93]), .CP(srdy), .Q(
        \input_weight_loc[2][13] ) );
  DFQD1 \input_weight_loc_reg[2][12]  ( .D(input_weight[92]), .CP(srdy), .Q(
        \input_weight_loc[2][12] ) );
  DFQD1 \input_weight_loc_reg[2][11]  ( .D(input_weight[91]), .CP(srdy), .Q(
        \input_weight_loc[2][11] ) );
  DFQD1 \input_weight_loc_reg[2][10]  ( .D(input_weight[90]), .CP(srdy), .Q(
        \input_weight_loc[2][10] ) );
  DFQD1 \input_weight_loc_reg[2][9]  ( .D(input_weight[89]), .CP(srdy), .Q(
        \input_weight_loc[2][9] ) );
  DFQD1 \input_weight_loc_reg[2][8]  ( .D(input_weight[88]), .CP(srdy), .Q(
        \input_weight_loc[2][8] ) );
  DFQD1 \input_weight_loc_reg[2][7]  ( .D(input_weight[87]), .CP(srdy), .Q(
        \input_weight_loc[2][7] ) );
  DFQD1 \input_weight_loc_reg[2][6]  ( .D(input_weight[86]), .CP(srdy), .Q(
        \input_weight_loc[2][6] ) );
  DFQD1 \input_weight_loc_reg[2][5]  ( .D(input_weight[85]), .CP(srdy), .Q(
        \input_weight_loc[2][5] ) );
  DFQD1 \input_weight_loc_reg[2][4]  ( .D(input_weight[84]), .CP(srdy), .Q(
        \input_weight_loc[2][4] ) );
  DFQD1 \input_weight_loc_reg[2][3]  ( .D(input_weight[83]), .CP(srdy), .Q(
        \input_weight_loc[2][3] ) );
  DFQD1 \input_weight_loc_reg[2][2]  ( .D(input_weight[82]), .CP(srdy), .Q(
        \input_weight_loc[2][2] ) );
  DFQD1 \input_weight_loc_reg[2][1]  ( .D(input_weight[81]), .CP(srdy), .Q(
        \input_weight_loc[2][1] ) );
  DFQD1 \input_weight_loc_reg[2][0]  ( .D(input_weight[80]), .CP(srdy), .Q(
        \input_weight_loc[2][0] ) );
  DFQD1 \input_weight_loc_reg[0][15]  ( .D(input_weight[127]), .CP(srdy), .Q(
        \input_weight_loc[0][15] ) );
  DFQD1 \input_weight_loc_reg[0][14]  ( .D(input_weight[126]), .CP(srdy), .Q(
        \input_weight_loc[0][14] ) );
  DFQD1 \input_weight_loc_reg[0][13]  ( .D(input_weight[125]), .CP(srdy), .Q(
        \input_weight_loc[0][13] ) );
  DFQD1 \input_weight_loc_reg[0][12]  ( .D(input_weight[124]), .CP(srdy), .Q(
        \input_weight_loc[0][12] ) );
  DFQD1 \input_weight_loc_reg[0][11]  ( .D(input_weight[123]), .CP(srdy), .Q(
        \input_weight_loc[0][11] ) );
  DFQD1 \input_weight_loc_reg[0][10]  ( .D(input_weight[122]), .CP(srdy), .Q(
        \input_weight_loc[0][10] ) );
  DFQD1 \input_weight_loc_reg[0][9]  ( .D(input_weight[121]), .CP(srdy), .Q(
        \input_weight_loc[0][9] ) );
  DFQD1 \input_weight_loc_reg[0][8]  ( .D(input_weight[120]), .CP(srdy), .Q(
        \input_weight_loc[0][8] ) );
  DFQD1 \input_weight_loc_reg[0][7]  ( .D(input_weight[119]), .CP(srdy), .Q(
        \input_weight_loc[0][7] ) );
  DFQD1 \input_weight_loc_reg[0][6]  ( .D(input_weight[118]), .CP(srdy), .Q(
        \input_weight_loc[0][6] ) );
  DFQD1 \input_weight_loc_reg[0][5]  ( .D(input_weight[117]), .CP(srdy), .Q(
        \input_weight_loc[0][5] ) );
  DFQD1 \input_weight_loc_reg[0][4]  ( .D(input_weight[116]), .CP(srdy), .Q(
        \input_weight_loc[0][4] ) );
  DFQD1 \input_weight_loc_reg[0][3]  ( .D(input_weight[115]), .CP(srdy), .Q(
        \input_weight_loc[0][3] ) );
  DFQD1 \input_weight_loc_reg[0][2]  ( .D(input_weight[114]), .CP(srdy), .Q(
        \input_weight_loc[0][2] ) );
  DFQD1 \input_weight_loc_reg[0][1]  ( .D(input_weight[113]), .CP(srdy), .Q(
        \input_weight_loc[0][1] ) );
  DFQD1 \input_weight_loc_reg[0][0]  ( .D(input_weight[112]), .CP(srdy), .Q(
        \input_weight_loc[0][0] ) );
  DFQD1 \input_value_loc_reg[7][15]  ( .D(input_value[15]), .CP(srdy), .Q(
        \input_value_loc[7][15] ) );
  DFQD1 \input_value_loc_reg[7][14]  ( .D(input_value[14]), .CP(srdy), .Q(
        \input_value_loc[7][14] ) );
  DFQD1 \input_value_loc_reg[7][13]  ( .D(input_value[13]), .CP(srdy), .Q(
        \input_value_loc[7][13] ) );
  DFQD1 \input_value_loc_reg[7][12]  ( .D(input_value[12]), .CP(srdy), .Q(
        \input_value_loc[7][12] ) );
  DFQD1 \input_value_loc_reg[7][11]  ( .D(input_value[11]), .CP(srdy), .Q(
        \input_value_loc[7][11] ) );
  DFQD1 \input_value_loc_reg[7][10]  ( .D(input_value[10]), .CP(srdy), .Q(
        \input_value_loc[7][10] ) );
  DFQD1 \input_value_loc_reg[7][9]  ( .D(input_value[9]), .CP(srdy), .Q(
        \input_value_loc[7][9] ) );
  DFQD1 \input_value_loc_reg[7][8]  ( .D(input_value[8]), .CP(srdy), .Q(
        \input_value_loc[7][8] ) );
  DFQD1 \input_value_loc_reg[7][7]  ( .D(input_value[7]), .CP(srdy), .Q(
        \input_value_loc[7][7] ) );
  DFQD1 \input_value_loc_reg[7][6]  ( .D(input_value[6]), .CP(srdy), .Q(
        \input_value_loc[7][6] ) );
  DFQD1 \input_value_loc_reg[7][5]  ( .D(input_value[5]), .CP(srdy), .Q(
        \input_value_loc[7][5] ) );
  DFQD1 \input_value_loc_reg[7][4]  ( .D(input_value[4]), .CP(srdy), .Q(
        \input_value_loc[7][4] ) );
  DFQD1 \input_value_loc_reg[7][3]  ( .D(input_value[3]), .CP(srdy), .Q(
        \input_value_loc[7][3] ) );
  DFQD1 \input_value_loc_reg[7][2]  ( .D(input_value[2]), .CP(srdy), .Q(
        \input_value_loc[7][2] ) );
  DFQD1 \input_value_loc_reg[7][1]  ( .D(input_value[1]), .CP(srdy), .Q(
        \input_value_loc[7][1] ) );
  DFQD1 \input_value_loc_reg[4][15]  ( .D(input_value[63]), .CP(srdy), .Q(
        \input_value_loc[4][15] ) );
  DFQD1 \input_value_loc_reg[4][14]  ( .D(input_value[62]), .CP(srdy), .Q(
        \input_value_loc[4][14] ) );
  DFQD1 \input_value_loc_reg[4][13]  ( .D(input_value[61]), .CP(srdy), .Q(
        \input_value_loc[4][13] ) );
  DFQD1 \input_value_loc_reg[4][12]  ( .D(input_value[60]), .CP(srdy), .Q(
        \input_value_loc[4][12] ) );
  DFQD1 \input_value_loc_reg[4][11]  ( .D(input_value[59]), .CP(srdy), .Q(
        \input_value_loc[4][11] ) );
  DFQD1 \input_value_loc_reg[4][10]  ( .D(input_value[58]), .CP(srdy), .Q(
        \input_value_loc[4][10] ) );
  DFQD1 \input_value_loc_reg[4][9]  ( .D(input_value[57]), .CP(srdy), .Q(
        \input_value_loc[4][9] ) );
  DFQD1 \input_value_loc_reg[4][8]  ( .D(input_value[56]), .CP(srdy), .Q(
        \input_value_loc[4][8] ) );
  DFQD1 \input_value_loc_reg[4][7]  ( .D(input_value[55]), .CP(srdy), .Q(
        \input_value_loc[4][7] ) );
  DFQD1 \input_value_loc_reg[4][6]  ( .D(input_value[54]), .CP(srdy), .Q(
        \input_value_loc[4][6] ) );
  DFQD1 \input_value_loc_reg[4][5]  ( .D(input_value[53]), .CP(srdy), .Q(
        \input_value_loc[4][5] ) );
  DFQD1 \input_value_loc_reg[4][4]  ( .D(input_value[52]), .CP(srdy), .Q(
        \input_value_loc[4][4] ) );
  DFQD1 \input_value_loc_reg[4][3]  ( .D(input_value[51]), .CP(srdy), .Q(
        \input_value_loc[4][3] ) );
  DFQD1 \input_value_loc_reg[4][2]  ( .D(input_value[50]), .CP(srdy), .Q(
        \input_value_loc[4][2] ) );
  DFQD1 \input_value_loc_reg[4][1]  ( .D(input_value[49]), .CP(srdy), .Q(
        \input_value_loc[4][1] ) );
  DFQD1 \input_value_loc_reg[4][0]  ( .D(input_value[48]), .CP(srdy), .Q(
        \input_value_loc[4][0] ) );
  DFQD1 \input_value_loc_reg[2][15]  ( .D(input_value[95]), .CP(srdy), .Q(
        \input_value_loc[2][15] ) );
  DFQD1 \input_value_loc_reg[2][14]  ( .D(input_value[94]), .CP(srdy), .Q(
        \input_value_loc[2][14] ) );
  DFQD1 \input_value_loc_reg[2][13]  ( .D(input_value[93]), .CP(srdy), .Q(
        \input_value_loc[2][13] ) );
  DFQD1 \input_value_loc_reg[2][12]  ( .D(input_value[92]), .CP(srdy), .Q(
        \input_value_loc[2][12] ) );
  DFQD1 \input_value_loc_reg[2][11]  ( .D(input_value[91]), .CP(srdy), .Q(
        \input_value_loc[2][11] ) );
  DFQD1 \input_value_loc_reg[2][10]  ( .D(input_value[90]), .CP(srdy), .Q(
        \input_value_loc[2][10] ) );
  DFQD1 \input_value_loc_reg[2][9]  ( .D(input_value[89]), .CP(srdy), .Q(
        \input_value_loc[2][9] ) );
  DFQD1 \input_value_loc_reg[2][8]  ( .D(input_value[88]), .CP(srdy), .Q(
        \input_value_loc[2][8] ) );
  DFQD1 \input_value_loc_reg[2][7]  ( .D(input_value[87]), .CP(srdy), .Q(
        \input_value_loc[2][7] ) );
  DFQD1 \input_value_loc_reg[2][6]  ( .D(input_value[86]), .CP(srdy), .Q(
        \input_value_loc[2][6] ) );
  DFQD1 \input_value_loc_reg[2][5]  ( .D(input_value[85]), .CP(srdy), .Q(
        \input_value_loc[2][5] ) );
  DFQD1 \input_value_loc_reg[2][4]  ( .D(input_value[84]), .CP(srdy), .Q(
        \input_value_loc[2][4] ) );
  DFQD1 \input_value_loc_reg[2][3]  ( .D(input_value[83]), .CP(srdy), .Q(
        \input_value_loc[2][3] ) );
  DFQD1 \input_value_loc_reg[2][2]  ( .D(input_value[82]), .CP(srdy), .Q(
        \input_value_loc[2][2] ) );
  DFQD1 \input_value_loc_reg[2][1]  ( .D(input_value[81]), .CP(srdy), .Q(
        \input_value_loc[2][1] ) );
  DFQD1 \input_value_loc_reg[2][0]  ( .D(input_value[80]), .CP(srdy), .Q(
        \input_value_loc[2][0] ) );
  DFQD1 \input_value_loc_reg[0][15]  ( .D(input_value[127]), .CP(srdy), .Q(
        \input_value_loc[0][15] ) );
  DFQD1 \input_value_loc_reg[0][14]  ( .D(input_value[126]), .CP(srdy), .Q(
        \input_value_loc[0][14] ) );
  DFQD1 \input_value_loc_reg[0][13]  ( .D(input_value[125]), .CP(srdy), .Q(
        \input_value_loc[0][13] ) );
  DFQD1 \input_value_loc_reg[0][12]  ( .D(input_value[124]), .CP(srdy), .Q(
        \input_value_loc[0][12] ) );
  DFQD1 \input_value_loc_reg[0][11]  ( .D(input_value[123]), .CP(srdy), .Q(
        \input_value_loc[0][11] ) );
  DFQD1 \input_value_loc_reg[0][10]  ( .D(input_value[122]), .CP(srdy), .Q(
        \input_value_loc[0][10] ) );
  DFQD1 \input_value_loc_reg[0][9]  ( .D(input_value[121]), .CP(srdy), .Q(
        \input_value_loc[0][9] ) );
  DFQD1 \input_value_loc_reg[0][8]  ( .D(input_value[120]), .CP(srdy), .Q(
        \input_value_loc[0][8] ) );
  DFQD1 \input_value_loc_reg[0][7]  ( .D(input_value[119]), .CP(srdy), .Q(
        \input_value_loc[0][7] ) );
  DFQD1 \input_value_loc_reg[0][6]  ( .D(input_value[118]), .CP(srdy), .Q(
        \input_value_loc[0][6] ) );
  DFQD1 \input_value_loc_reg[0][5]  ( .D(input_value[117]), .CP(srdy), .Q(
        \input_value_loc[0][5] ) );
  DFQD1 \input_value_loc_reg[0][4]  ( .D(input_value[116]), .CP(srdy), .Q(
        \input_value_loc[0][4] ) );
  DFQD1 \input_value_loc_reg[0][3]  ( .D(input_value[115]), .CP(srdy), .Q(
        \input_value_loc[0][3] ) );
  DFQD1 \input_value_loc_reg[0][2]  ( .D(input_value[114]), .CP(srdy), .Q(
        \input_value_loc[0][2] ) );
  DFQD1 \input_value_loc_reg[0][1]  ( .D(input_value[113]), .CP(srdy), .Q(
        \input_value_loc[0][1] ) );
  DFQD1 \input_value_loc_reg[0][0]  ( .D(input_value[112]), .CP(srdy), .Q(
        \input_value_loc[0][0] ) );
  DFQD1 \input_weight_loc_reg[5][15]  ( .D(input_weight[47]), .CP(srdy), .Q(
        \input_weight_loc[5][15] ) );
  DFQD1 \input_weight_loc_reg[5][14]  ( .D(input_weight[46]), .CP(srdy), .Q(
        \input_weight_loc[5][14] ) );
  DFQD1 \input_weight_loc_reg[5][13]  ( .D(input_weight[45]), .CP(srdy), .Q(
        \input_weight_loc[5][13] ) );
  DFQD1 \input_weight_loc_reg[5][12]  ( .D(input_weight[44]), .CP(srdy), .Q(
        \input_weight_loc[5][12] ) );
  DFQD1 \input_weight_loc_reg[5][11]  ( .D(input_weight[43]), .CP(srdy), .Q(
        \input_weight_loc[5][11] ) );
  DFQD1 \input_weight_loc_reg[5][10]  ( .D(input_weight[42]), .CP(srdy), .Q(
        \input_weight_loc[5][10] ) );
  DFQD1 \input_weight_loc_reg[5][9]  ( .D(input_weight[41]), .CP(srdy), .Q(
        \input_weight_loc[5][9] ) );
  DFQD1 \input_weight_loc_reg[5][8]  ( .D(input_weight[40]), .CP(srdy), .Q(
        \input_weight_loc[5][8] ) );
  DFQD1 \input_weight_loc_reg[5][7]  ( .D(input_weight[39]), .CP(srdy), .Q(
        \input_weight_loc[5][7] ) );
  DFQD1 \input_weight_loc_reg[5][6]  ( .D(input_weight[38]), .CP(srdy), .Q(
        \input_weight_loc[5][6] ) );
  DFQD1 \input_weight_loc_reg[5][5]  ( .D(input_weight[37]), .CP(srdy), .Q(
        \input_weight_loc[5][5] ) );
  DFQD1 \input_weight_loc_reg[5][4]  ( .D(input_weight[36]), .CP(srdy), .Q(
        \input_weight_loc[5][4] ) );
  DFQD1 \input_weight_loc_reg[5][3]  ( .D(input_weight[35]), .CP(srdy), .Q(
        \input_weight_loc[5][3] ) );
  DFQD1 \input_weight_loc_reg[5][2]  ( .D(input_weight[34]), .CP(srdy), .Q(
        \input_weight_loc[5][2] ) );
  DFQD1 \input_weight_loc_reg[5][1]  ( .D(input_weight[33]), .CP(srdy), .Q(
        \input_weight_loc[5][1] ) );
  DFQD1 \input_weight_loc_reg[5][0]  ( .D(input_weight[32]), .CP(srdy), .Q(
        \input_weight_loc[5][0] ) );
  DFQD1 \input_value_loc_reg[5][0]  ( .D(input_value[32]), .CP(srdy), .Q(
        \input_value_loc[5][0] ) );
  DFQD1 \output_value_loc_reg[0]  ( .D(fma_z[0]), .CP(\*Logic1* ), .Q(
        output_value_loc[0]) );
  DFQD1 \output_value_loc_reg[1]  ( .D(fma_z[1]), .CP(\*Logic1* ), .Q(
        output_value_loc[1]) );
  DFQD1 \output_value_loc_reg[2]  ( .D(fma_z[2]), .CP(\*Logic1* ), .Q(
        output_value_loc[2]) );
  DFQD1 \output_value_loc_reg[3]  ( .D(fma_z[3]), .CP(\*Logic1* ), .Q(
        output_value_loc[3]) );
  DFQD1 \output_value_loc_reg[4]  ( .D(fma_z[4]), .CP(\*Logic1* ), .Q(
        output_value_loc[4]) );
  DFQD1 \output_value_loc_reg[5]  ( .D(fma_z[5]), .CP(\*Logic1* ), .Q(
        output_value_loc[5]) );
  DFQD1 \output_value_loc_reg[6]  ( .D(fma_z[6]), .CP(\*Logic1* ), .Q(
        output_value_loc[6]) );
  DFQD1 \output_value_loc_reg[7]  ( .D(fma_z[7]), .CP(\*Logic1* ), .Q(
        output_value_loc[7]) );
  DFQD1 \output_value_loc_reg[8]  ( .D(fma_z[8]), .CP(\*Logic1* ), .Q(
        output_value_loc[8]) );
  DFQD1 \output_value_loc_reg[9]  ( .D(fma_z[9]), .CP(\*Logic1* ), .Q(
        output_value_loc[9]) );
  DFQD1 \output_value_loc_reg[10]  ( .D(fma_z[10]), .CP(\*Logic1* ), .Q(
        output_value_loc[10]) );
  DFQD1 \output_value_loc_reg[11]  ( .D(fma_z[11]), .CP(\*Logic1* ), .Q(
        output_value_loc[11]) );
  DFQD1 \output_value_loc_reg[12]  ( .D(fma_z[12]), .CP(\*Logic1* ), .Q(
        output_value_loc[12]) );
  DFQD1 \output_value_loc_reg[13]  ( .D(fma_z[13]), .CP(\*Logic1* ), .Q(
        output_value_loc[13]) );
  DFQD1 \output_value_loc_reg[14]  ( .D(fma_z[14]), .CP(\*Logic1* ), .Q(
        output_value_loc[14]) );
  DFQD1 \output_value_loc_reg[15]  ( .D(n1), .CP(\*Logic1* ), .Q(
        output_value_loc[15]) );
  DFQD1 \input_weight_loc_reg[7][15]  ( .D(input_weight[15]), .CP(srdy), .Q(
        \input_weight_loc[7][15] ) );
  DFQD1 \input_weight_loc_reg[7][14]  ( .D(input_weight[14]), .CP(srdy), .Q(
        \input_weight_loc[7][14] ) );
  DFQD1 \input_weight_loc_reg[7][13]  ( .D(input_weight[13]), .CP(srdy), .Q(
        \input_weight_loc[7][13] ) );
  DFQD1 \input_weight_loc_reg[7][12]  ( .D(input_weight[12]), .CP(srdy), .Q(
        \input_weight_loc[7][12] ) );
  DFQD1 \input_weight_loc_reg[7][11]  ( .D(input_weight[11]), .CP(srdy), .Q(
        \input_weight_loc[7][11] ) );
  DFQD1 \input_weight_loc_reg[7][10]  ( .D(input_weight[10]), .CP(srdy), .Q(
        \input_weight_loc[7][10] ) );
  DFQD1 \input_weight_loc_reg[7][9]  ( .D(input_weight[9]), .CP(srdy), .Q(
        \input_weight_loc[7][9] ) );
  DFQD1 \input_weight_loc_reg[7][8]  ( .D(input_weight[8]), .CP(srdy), .Q(
        \input_weight_loc[7][8] ) );
  DFQD1 \input_weight_loc_reg[7][7]  ( .D(input_weight[7]), .CP(srdy), .Q(
        \input_weight_loc[7][7] ) );
  DFQD1 \input_weight_loc_reg[7][6]  ( .D(input_weight[6]), .CP(srdy), .Q(
        \input_weight_loc[7][6] ) );
  DFQD1 \input_weight_loc_reg[7][5]  ( .D(input_weight[5]), .CP(srdy), .Q(
        \input_weight_loc[7][5] ) );
  DFQD1 \input_weight_loc_reg[7][4]  ( .D(input_weight[4]), .CP(srdy), .Q(
        \input_weight_loc[7][4] ) );
  DFQD1 \input_weight_loc_reg[7][3]  ( .D(input_weight[3]), .CP(srdy), .Q(
        \input_weight_loc[7][3] ) );
  DFQD1 \input_weight_loc_reg[7][2]  ( .D(input_weight[2]), .CP(srdy), .Q(
        \input_weight_loc[7][2] ) );
  DFQD1 \input_weight_loc_reg[7][1]  ( .D(input_weight[1]), .CP(srdy), .Q(
        \input_weight_loc[7][1] ) );
  DFQD1 \input_weight_loc_reg[7][0]  ( .D(input_weight[0]), .CP(srdy), .Q(
        \input_weight_loc[7][0] ) );
  DFQD1 \input_value_loc_reg[7][0]  ( .D(input_value[0]), .CP(srdy), .Q(
        \input_value_loc[7][0] ) );
  DFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .CP(\*Logic1* ), .Q(
        cur_state[2]) );
  DFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .CP(\*Logic1* ), .Q(
        cur_state[3]) );
  DFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .CP(\*Logic1* ), .Q(
        cur_state[1]) );
  DFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .CP(\*Logic1* ), .Q(
        cur_state[0]) );
  TIEL U3 ( .ZN(n1) );
  INR2XD0 U4 ( .A1(n57), .B1(n10), .ZN(n21) );
  IND4D1 U5 ( .A1(n3), .B1(n7), .B2(n12), .B3(n56), .ZN(N90) );
  NR4D1 U6 ( .A1(n4), .A2(cur_state[0]), .A3(cur_state[1]), .A4(cur_state[3]), 
        .ZN(n20) );
  TIEH U7 ( .Z(\*Logic1* ) );
  OR2D0 U8 ( .A1(n2), .A2(n3), .Z(nxt_state[3]) );
  OAI211D0 U9 ( .A1(n4), .A2(n5), .B(n6), .C(n7), .ZN(nxt_state[2]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n5) );
  OAI211D0 U11 ( .A1(cur_state[1]), .A2(n10), .B(n6), .C(n11), .ZN(
        nxt_state[1]) );
  CKND0 U12 ( .I(n12), .ZN(nxt_state[0]) );
  ND4D0 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(N99) );
  AOI22D0 U14 ( .A1(\input_value_loc[7][8] ), .A2(n2), .B1(
        \input_value_loc[5][8] ), .B2(n17), .ZN(n16) );
  AOI22D0 U15 ( .A1(\input_value_loc[4][8] ), .A2(n18), .B1(
        \input_value_loc[6][8] ), .B2(n3), .ZN(n15) );
  AOI22D0 U16 ( .A1(\input_value_loc[2][8] ), .A2(n19), .B1(
        \input_value_loc[3][8] ), .B2(n20), .ZN(n14) );
  AOI22D0 U17 ( .A1(\input_value_loc[0][8] ), .A2(n21), .B1(
        \input_value_loc[1][8] ), .B2(n22), .ZN(n13) );
  ND4D0 U18 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(N98) );
  AOI22D0 U19 ( .A1(\input_value_loc[7][7] ), .A2(n2), .B1(
        \input_value_loc[5][7] ), .B2(n17), .ZN(n26) );
  AOI22D0 U20 ( .A1(\input_value_loc[4][7] ), .A2(n18), .B1(
        \input_value_loc[6][7] ), .B2(n3), .ZN(n25) );
  AOI22D0 U21 ( .A1(\input_value_loc[2][7] ), .A2(n19), .B1(
        \input_value_loc[3][7] ), .B2(n20), .ZN(n24) );
  AOI22D0 U22 ( .A1(\input_value_loc[0][7] ), .A2(n21), .B1(
        \input_value_loc[1][7] ), .B2(n22), .ZN(n23) );
  ND4D0 U23 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(N97) );
  AOI22D0 U24 ( .A1(\input_value_loc[7][6] ), .A2(n2), .B1(
        \input_value_loc[5][6] ), .B2(n17), .ZN(n30) );
  AOI22D0 U25 ( .A1(\input_value_loc[4][6] ), .A2(n18), .B1(
        \input_value_loc[6][6] ), .B2(n3), .ZN(n29) );
  AOI22D0 U26 ( .A1(\input_value_loc[2][6] ), .A2(n19), .B1(
        \input_value_loc[3][6] ), .B2(n20), .ZN(n28) );
  AOI22D0 U27 ( .A1(\input_value_loc[0][6] ), .A2(n21), .B1(
        \input_value_loc[1][6] ), .B2(n22), .ZN(n27) );
  ND4D0 U28 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(N96) );
  AOI22D0 U29 ( .A1(\input_value_loc[7][5] ), .A2(n2), .B1(
        \input_value_loc[5][5] ), .B2(n17), .ZN(n34) );
  AOI22D0 U30 ( .A1(\input_value_loc[4][5] ), .A2(n18), .B1(
        \input_value_loc[6][5] ), .B2(n3), .ZN(n33) );
  AOI22D0 U31 ( .A1(\input_value_loc[2][5] ), .A2(n19), .B1(
        \input_value_loc[3][5] ), .B2(n20), .ZN(n32) );
  AOI22D0 U32 ( .A1(\input_value_loc[0][5] ), .A2(n21), .B1(
        \input_value_loc[1][5] ), .B2(n22), .ZN(n31) );
  ND4D0 U33 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(N95) );
  AOI22D0 U34 ( .A1(\input_value_loc[7][4] ), .A2(n2), .B1(
        \input_value_loc[5][4] ), .B2(n17), .ZN(n38) );
  AOI22D0 U35 ( .A1(\input_value_loc[4][4] ), .A2(n18), .B1(
        \input_value_loc[6][4] ), .B2(n3), .ZN(n37) );
  AOI22D0 U36 ( .A1(\input_value_loc[2][4] ), .A2(n19), .B1(
        \input_value_loc[3][4] ), .B2(n20), .ZN(n36) );
  AOI22D0 U37 ( .A1(\input_value_loc[0][4] ), .A2(n21), .B1(
        \input_value_loc[1][4] ), .B2(n22), .ZN(n35) );
  ND4D0 U38 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(N94) );
  AOI22D0 U39 ( .A1(\input_value_loc[7][3] ), .A2(n2), .B1(
        \input_value_loc[5][3] ), .B2(n17), .ZN(n42) );
  AOI22D0 U40 ( .A1(\input_value_loc[4][3] ), .A2(n18), .B1(
        \input_value_loc[6][3] ), .B2(n3), .ZN(n41) );
  AOI22D0 U41 ( .A1(\input_value_loc[2][3] ), .A2(n19), .B1(
        \input_value_loc[3][3] ), .B2(n20), .ZN(n40) );
  AOI22D0 U42 ( .A1(\input_value_loc[0][3] ), .A2(n21), .B1(
        \input_value_loc[1][3] ), .B2(n22), .ZN(n39) );
  ND4D0 U43 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(N93) );
  AOI22D0 U44 ( .A1(\input_value_loc[7][2] ), .A2(n2), .B1(
        \input_value_loc[5][2] ), .B2(n17), .ZN(n46) );
  AOI22D0 U45 ( .A1(\input_value_loc[4][2] ), .A2(n18), .B1(
        \input_value_loc[6][2] ), .B2(n3), .ZN(n45) );
  AOI22D0 U46 ( .A1(\input_value_loc[2][2] ), .A2(n19), .B1(
        \input_value_loc[3][2] ), .B2(n20), .ZN(n44) );
  AOI22D0 U47 ( .A1(\input_value_loc[0][2] ), .A2(n21), .B1(
        \input_value_loc[1][2] ), .B2(n22), .ZN(n43) );
  ND4D0 U48 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(N92) );
  AOI22D0 U49 ( .A1(\input_value_loc[7][1] ), .A2(n2), .B1(
        \input_value_loc[5][1] ), .B2(n17), .ZN(n50) );
  AOI22D0 U50 ( .A1(\input_value_loc[4][1] ), .A2(n18), .B1(
        \input_value_loc[6][1] ), .B2(n3), .ZN(n49) );
  AOI22D0 U51 ( .A1(\input_value_loc[2][1] ), .A2(n19), .B1(
        \input_value_loc[3][1] ), .B2(n20), .ZN(n48) );
  AOI22D0 U52 ( .A1(\input_value_loc[0][1] ), .A2(n21), .B1(
        \input_value_loc[1][1] ), .B2(n22), .ZN(n47) );
  ND4D0 U53 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(N91) );
  AOI221D0 U54 ( .A1(\input_value_loc[5][0] ), .A2(n17), .B1(
        \input_value_loc[7][0] ), .B2(n2), .C(n55), .ZN(n54) );
  AOI22D0 U55 ( .A1(\input_value_loc[4][0] ), .A2(n18), .B1(
        \input_value_loc[6][0] ), .B2(n3), .ZN(n53) );
  AOI22D0 U56 ( .A1(\input_value_loc[2][0] ), .A2(n19), .B1(
        \input_value_loc[3][0] ), .B2(n20), .ZN(n52) );
  AOI22D0 U57 ( .A1(\input_value_loc[0][0] ), .A2(n21), .B1(
        \input_value_loc[1][0] ), .B2(n22), .ZN(n51) );
  NR2D0 U58 ( .A1(n18), .A2(n57), .ZN(n56) );
  NR4D0 U59 ( .A1(n20), .A2(n2), .A3(n17), .A4(n22), .ZN(n12) );
  CKND0 U60 ( .I(n19), .ZN(n7) );
  ND4D0 U61 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(N122) );
  AOI222D0 U62 ( .A1(\input_weight_loc[5][15] ), .A2(n17), .B1(
        output_value_loc[15]), .B2(n55), .C1(\input_weight_loc[7][15] ), .C2(
        n2), .ZN(n61) );
  AOI22D0 U63 ( .A1(\input_weight_loc[4][15] ), .A2(n18), .B1(
        \input_weight_loc[6][15] ), .B2(n3), .ZN(n60) );
  AOI22D0 U64 ( .A1(\input_weight_loc[2][15] ), .A2(n19), .B1(
        \input_weight_loc[3][15] ), .B2(n20), .ZN(n59) );
  AOI22D0 U65 ( .A1(\input_weight_loc[0][15] ), .A2(n21), .B1(
        \input_weight_loc[1][15] ), .B2(n22), .ZN(n58) );
  ND4D0 U66 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(N121) );
  AOI222D0 U67 ( .A1(\input_weight_loc[5][14] ), .A2(n17), .B1(
        output_value_loc[14]), .B2(n55), .C1(\input_weight_loc[7][14] ), .C2(
        n2), .ZN(n65) );
  AOI22D0 U68 ( .A1(\input_weight_loc[4][14] ), .A2(n18), .B1(
        \input_weight_loc[6][14] ), .B2(n3), .ZN(n64) );
  AOI22D0 U69 ( .A1(\input_weight_loc[2][14] ), .A2(n19), .B1(
        \input_weight_loc[3][14] ), .B2(n20), .ZN(n63) );
  AOI22D0 U70 ( .A1(\input_weight_loc[0][14] ), .A2(n21), .B1(
        \input_weight_loc[1][14] ), .B2(n22), .ZN(n62) );
  ND4D0 U71 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(N120) );
  AOI222D0 U72 ( .A1(\input_weight_loc[5][13] ), .A2(n17), .B1(
        output_value_loc[13]), .B2(n55), .C1(\input_weight_loc[7][13] ), .C2(
        n2), .ZN(n69) );
  AOI22D0 U73 ( .A1(\input_weight_loc[4][13] ), .A2(n18), .B1(
        \input_weight_loc[6][13] ), .B2(n3), .ZN(n68) );
  AOI22D0 U74 ( .A1(\input_weight_loc[2][13] ), .A2(n19), .B1(
        \input_weight_loc[3][13] ), .B2(n20), .ZN(n67) );
  AOI22D0 U75 ( .A1(\input_weight_loc[0][13] ), .A2(n21), .B1(
        \input_weight_loc[1][13] ), .B2(n22), .ZN(n66) );
  ND4D0 U76 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(N119) );
  AOI222D0 U77 ( .A1(\input_weight_loc[5][12] ), .A2(n17), .B1(
        output_value_loc[12]), .B2(n55), .C1(\input_weight_loc[7][12] ), .C2(
        n2), .ZN(n73) );
  AOI22D0 U78 ( .A1(\input_weight_loc[4][12] ), .A2(n18), .B1(
        \input_weight_loc[6][12] ), .B2(n3), .ZN(n72) );
  AOI22D0 U79 ( .A1(\input_weight_loc[2][12] ), .A2(n19), .B1(
        \input_weight_loc[3][12] ), .B2(n20), .ZN(n71) );
  AOI22D0 U80 ( .A1(\input_weight_loc[0][12] ), .A2(n21), .B1(
        \input_weight_loc[1][12] ), .B2(n22), .ZN(n70) );
  ND4D0 U81 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(N118) );
  AOI222D0 U82 ( .A1(\input_weight_loc[5][11] ), .A2(n17), .B1(
        output_value_loc[11]), .B2(n55), .C1(\input_weight_loc[7][11] ), .C2(
        n2), .ZN(n77) );
  AOI22D0 U83 ( .A1(\input_weight_loc[4][11] ), .A2(n18), .B1(
        \input_weight_loc[6][11] ), .B2(n3), .ZN(n76) );
  AOI22D0 U84 ( .A1(\input_weight_loc[2][11] ), .A2(n19), .B1(
        \input_weight_loc[3][11] ), .B2(n20), .ZN(n75) );
  AOI22D0 U85 ( .A1(\input_weight_loc[0][11] ), .A2(n21), .B1(
        \input_weight_loc[1][11] ), .B2(n22), .ZN(n74) );
  ND4D0 U86 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(N117) );
  AOI222D0 U87 ( .A1(\input_weight_loc[5][10] ), .A2(n17), .B1(
        output_value_loc[10]), .B2(n55), .C1(\input_weight_loc[7][10] ), .C2(
        n2), .ZN(n81) );
  AOI22D0 U88 ( .A1(\input_weight_loc[4][10] ), .A2(n18), .B1(
        \input_weight_loc[6][10] ), .B2(n3), .ZN(n80) );
  AOI22D0 U89 ( .A1(\input_weight_loc[2][10] ), .A2(n19), .B1(
        \input_weight_loc[3][10] ), .B2(n20), .ZN(n79) );
  AOI22D0 U90 ( .A1(\input_weight_loc[0][10] ), .A2(n21), .B1(
        \input_weight_loc[1][10] ), .B2(n22), .ZN(n78) );
  ND4D0 U91 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(N116) );
  AOI222D0 U92 ( .A1(\input_weight_loc[5][9] ), .A2(n17), .B1(
        output_value_loc[9]), .B2(n55), .C1(\input_weight_loc[7][9] ), .C2(n2), 
        .ZN(n85) );
  AOI22D0 U93 ( .A1(\input_weight_loc[4][9] ), .A2(n18), .B1(
        \input_weight_loc[6][9] ), .B2(n3), .ZN(n84) );
  AOI22D0 U94 ( .A1(\input_weight_loc[2][9] ), .A2(n19), .B1(
        \input_weight_loc[3][9] ), .B2(n20), .ZN(n83) );
  AOI22D0 U95 ( .A1(\input_weight_loc[0][9] ), .A2(n21), .B1(
        \input_weight_loc[1][9] ), .B2(n22), .ZN(n82) );
  ND4D0 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(N115) );
  AOI222D0 U97 ( .A1(\input_weight_loc[5][8] ), .A2(n17), .B1(
        output_value_loc[8]), .B2(n55), .C1(\input_weight_loc[7][8] ), .C2(n2), 
        .ZN(n89) );
  AOI22D0 U98 ( .A1(\input_weight_loc[4][8] ), .A2(n18), .B1(
        \input_weight_loc[6][8] ), .B2(n3), .ZN(n88) );
  AOI22D0 U99 ( .A1(\input_weight_loc[2][8] ), .A2(n19), .B1(
        \input_weight_loc[3][8] ), .B2(n20), .ZN(n87) );
  AOI22D0 U100 ( .A1(\input_weight_loc[0][8] ), .A2(n21), .B1(
        \input_weight_loc[1][8] ), .B2(n22), .ZN(n86) );
  ND4D0 U101 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(N114) );
  AOI222D0 U102 ( .A1(\input_weight_loc[5][7] ), .A2(n17), .B1(
        output_value_loc[7]), .B2(n55), .C1(\input_weight_loc[7][7] ), .C2(n2), 
        .ZN(n93) );
  AOI22D0 U103 ( .A1(\input_weight_loc[4][7] ), .A2(n18), .B1(
        \input_weight_loc[6][7] ), .B2(n3), .ZN(n92) );
  AOI22D0 U104 ( .A1(\input_weight_loc[2][7] ), .A2(n19), .B1(
        \input_weight_loc[3][7] ), .B2(n20), .ZN(n91) );
  AOI22D0 U105 ( .A1(\input_weight_loc[0][7] ), .A2(n21), .B1(
        \input_weight_loc[1][7] ), .B2(n22), .ZN(n90) );
  ND4D0 U106 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(N113) );
  AOI222D0 U107 ( .A1(\input_weight_loc[5][6] ), .A2(n17), .B1(
        output_value_loc[6]), .B2(n55), .C1(\input_weight_loc[7][6] ), .C2(n2), 
        .ZN(n97) );
  AOI22D0 U108 ( .A1(\input_weight_loc[4][6] ), .A2(n18), .B1(
        \input_weight_loc[6][6] ), .B2(n3), .ZN(n96) );
  AOI22D0 U109 ( .A1(\input_weight_loc[2][6] ), .A2(n19), .B1(
        \input_weight_loc[3][6] ), .B2(n20), .ZN(n95) );
  AOI22D0 U110 ( .A1(\input_weight_loc[0][6] ), .A2(n21), .B1(
        \input_weight_loc[1][6] ), .B2(n22), .ZN(n94) );
  ND4D0 U111 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(N112) );
  AOI222D0 U112 ( .A1(\input_weight_loc[5][5] ), .A2(n17), .B1(
        output_value_loc[5]), .B2(n55), .C1(\input_weight_loc[7][5] ), .C2(n2), 
        .ZN(n101) );
  AOI22D0 U113 ( .A1(\input_weight_loc[4][5] ), .A2(n18), .B1(
        \input_weight_loc[6][5] ), .B2(n3), .ZN(n100) );
  AOI22D0 U114 ( .A1(\input_weight_loc[2][5] ), .A2(n19), .B1(
        \input_weight_loc[3][5] ), .B2(n20), .ZN(n99) );
  AOI22D0 U115 ( .A1(\input_weight_loc[0][5] ), .A2(n21), .B1(
        \input_weight_loc[1][5] ), .B2(n22), .ZN(n98) );
  ND4D0 U116 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(N111) );
  AOI222D0 U117 ( .A1(\input_weight_loc[5][4] ), .A2(n17), .B1(
        output_value_loc[4]), .B2(n55), .C1(\input_weight_loc[7][4] ), .C2(n2), 
        .ZN(n105) );
  AOI22D0 U118 ( .A1(\input_weight_loc[4][4] ), .A2(n18), .B1(
        \input_weight_loc[6][4] ), .B2(n3), .ZN(n104) );
  AOI22D0 U119 ( .A1(\input_weight_loc[2][4] ), .A2(n19), .B1(
        \input_weight_loc[3][4] ), .B2(n20), .ZN(n103) );
  AOI22D0 U120 ( .A1(\input_weight_loc[0][4] ), .A2(n21), .B1(
        \input_weight_loc[1][4] ), .B2(n22), .ZN(n102) );
  ND4D0 U121 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(N110) );
  AOI222D0 U122 ( .A1(\input_weight_loc[5][3] ), .A2(n17), .B1(
        output_value_loc[3]), .B2(n55), .C1(\input_weight_loc[7][3] ), .C2(n2), 
        .ZN(n109) );
  AOI22D0 U123 ( .A1(\input_weight_loc[4][3] ), .A2(n18), .B1(
        \input_weight_loc[6][3] ), .B2(n3), .ZN(n108) );
  AOI22D0 U124 ( .A1(\input_weight_loc[2][3] ), .A2(n19), .B1(
        \input_weight_loc[3][3] ), .B2(n20), .ZN(n107) );
  AOI22D0 U125 ( .A1(\input_weight_loc[0][3] ), .A2(n21), .B1(
        \input_weight_loc[1][3] ), .B2(n22), .ZN(n106) );
  ND4D0 U126 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(N109) );
  AOI222D0 U127 ( .A1(\input_weight_loc[5][2] ), .A2(n17), .B1(
        output_value_loc[2]), .B2(n55), .C1(\input_weight_loc[7][2] ), .C2(n2), 
        .ZN(n113) );
  AOI22D0 U128 ( .A1(\input_weight_loc[4][2] ), .A2(n18), .B1(
        \input_weight_loc[6][2] ), .B2(n3), .ZN(n112) );
  AOI22D0 U129 ( .A1(\input_weight_loc[2][2] ), .A2(n19), .B1(
        \input_weight_loc[3][2] ), .B2(n20), .ZN(n111) );
  AOI22D0 U130 ( .A1(\input_weight_loc[0][2] ), .A2(n21), .B1(
        \input_weight_loc[1][2] ), .B2(n22), .ZN(n110) );
  ND4D0 U131 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .ZN(N108) );
  AOI222D0 U132 ( .A1(\input_weight_loc[5][1] ), .A2(n17), .B1(
        output_value_loc[1]), .B2(n55), .C1(\input_weight_loc[7][1] ), .C2(n2), 
        .ZN(n117) );
  AOI22D0 U133 ( .A1(\input_weight_loc[4][1] ), .A2(n18), .B1(
        \input_weight_loc[6][1] ), .B2(n3), .ZN(n116) );
  AOI22D0 U134 ( .A1(\input_weight_loc[2][1] ), .A2(n19), .B1(
        \input_weight_loc[3][1] ), .B2(n20), .ZN(n115) );
  AOI22D0 U135 ( .A1(\input_weight_loc[0][1] ), .A2(n21), .B1(
        \input_weight_loc[1][1] ), .B2(n22), .ZN(n114) );
  ND4D0 U136 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(N107) );
  AOI222D0 U137 ( .A1(\input_weight_loc[5][0] ), .A2(n17), .B1(
        output_value_loc[0]), .B2(n55), .C1(\input_weight_loc[7][0] ), .C2(n2), 
        .ZN(n121) );
  AN3D0 U138 ( .A1(cur_state[3]), .A2(n57), .A3(cur_state[0]), .Z(n55) );
  AOI22D0 U139 ( .A1(\input_weight_loc[4][0] ), .A2(n18), .B1(
        \input_weight_loc[6][0] ), .B2(n3), .ZN(n120) );
  AOI22D0 U140 ( .A1(\input_weight_loc[2][0] ), .A2(n19), .B1(
        \input_weight_loc[3][0] ), .B2(n20), .ZN(n119) );
  AOI22D0 U141 ( .A1(\input_weight_loc[0][0] ), .A2(n21), .B1(
        \input_weight_loc[1][0] ), .B2(n22), .ZN(n118) );
  ND4D0 U142 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(N106) );
  AOI22D0 U143 ( .A1(\input_value_loc[7][15] ), .A2(n2), .B1(
        \input_value_loc[5][15] ), .B2(n17), .ZN(n125) );
  AOI22D0 U144 ( .A1(\input_value_loc[4][15] ), .A2(n18), .B1(
        \input_value_loc[6][15] ), .B2(n3), .ZN(n124) );
  AOI22D0 U145 ( .A1(\input_value_loc[2][15] ), .A2(n19), .B1(
        \input_value_loc[3][15] ), .B2(n20), .ZN(n123) );
  AOI22D0 U146 ( .A1(\input_value_loc[0][15] ), .A2(n21), .B1(
        \input_value_loc[1][15] ), .B2(n22), .ZN(n122) );
  ND4D0 U147 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(N105) );
  AOI22D0 U148 ( .A1(\input_value_loc[7][14] ), .A2(n2), .B1(
        \input_value_loc[5][14] ), .B2(n17), .ZN(n129) );
  AOI22D0 U149 ( .A1(\input_value_loc[4][14] ), .A2(n18), .B1(
        \input_value_loc[6][14] ), .B2(n3), .ZN(n128) );
  AOI22D0 U150 ( .A1(\input_value_loc[2][14] ), .A2(n19), .B1(
        \input_value_loc[3][14] ), .B2(n20), .ZN(n127) );
  AOI22D0 U151 ( .A1(\input_value_loc[0][14] ), .A2(n21), .B1(
        \input_value_loc[1][14] ), .B2(n22), .ZN(n126) );
  ND4D0 U152 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(N104) );
  AOI22D0 U153 ( .A1(\input_value_loc[7][13] ), .A2(n2), .B1(
        \input_value_loc[5][13] ), .B2(n17), .ZN(n133) );
  AOI22D0 U154 ( .A1(\input_value_loc[4][13] ), .A2(n18), .B1(
        \input_value_loc[6][13] ), .B2(n3), .ZN(n132) );
  AOI22D0 U155 ( .A1(\input_value_loc[2][13] ), .A2(n19), .B1(
        \input_value_loc[3][13] ), .B2(n20), .ZN(n131) );
  AOI22D0 U156 ( .A1(\input_value_loc[0][13] ), .A2(n21), .B1(
        \input_value_loc[1][13] ), .B2(n22), .ZN(n130) );
  ND4D0 U157 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(N103) );
  AOI22D0 U158 ( .A1(\input_value_loc[7][12] ), .A2(n2), .B1(
        \input_value_loc[5][12] ), .B2(n17), .ZN(n137) );
  AOI22D0 U159 ( .A1(\input_value_loc[4][12] ), .A2(n18), .B1(
        \input_value_loc[6][12] ), .B2(n3), .ZN(n136) );
  AOI22D0 U160 ( .A1(\input_value_loc[2][12] ), .A2(n19), .B1(
        \input_value_loc[3][12] ), .B2(n20), .ZN(n135) );
  AOI22D0 U161 ( .A1(\input_value_loc[0][12] ), .A2(n21), .B1(
        \input_value_loc[1][12] ), .B2(n22), .ZN(n134) );
  ND4D0 U162 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(N102) );
  AOI22D0 U163 ( .A1(\input_value_loc[7][11] ), .A2(n2), .B1(
        \input_value_loc[5][11] ), .B2(n17), .ZN(n141) );
  AOI22D0 U164 ( .A1(\input_value_loc[4][11] ), .A2(n18), .B1(
        \input_value_loc[6][11] ), .B2(n3), .ZN(n140) );
  AOI22D0 U165 ( .A1(\input_value_loc[2][11] ), .A2(n19), .B1(
        \input_value_loc[3][11] ), .B2(n20), .ZN(n139) );
  AOI22D0 U166 ( .A1(\input_value_loc[0][11] ), .A2(n21), .B1(
        \input_value_loc[1][11] ), .B2(n22), .ZN(n138) );
  ND4D0 U167 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(N101) );
  AOI22D0 U168 ( .A1(\input_value_loc[7][10] ), .A2(n2), .B1(
        \input_value_loc[5][10] ), .B2(n17), .ZN(n145) );
  AOI22D0 U169 ( .A1(\input_value_loc[4][10] ), .A2(n18), .B1(
        \input_value_loc[6][10] ), .B2(n3), .ZN(n144) );
  AOI22D0 U170 ( .A1(\input_value_loc[2][10] ), .A2(n19), .B1(
        \input_value_loc[3][10] ), .B2(n20), .ZN(n143) );
  AOI22D0 U171 ( .A1(\input_value_loc[0][10] ), .A2(n21), .B1(
        \input_value_loc[1][10] ), .B2(n22), .ZN(n142) );
  ND4D0 U172 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(N100) );
  AOI22D0 U173 ( .A1(\input_value_loc[7][9] ), .A2(n2), .B1(
        \input_value_loc[5][9] ), .B2(n17), .ZN(n149) );
  CKND0 U174 ( .I(n6), .ZN(n17) );
  CKND2D0 U175 ( .A1(n150), .A2(cur_state[2]), .ZN(n6) );
  INR3D0 U176 ( .A1(n57), .B1(cur_state[0]), .B2(n9), .ZN(n2) );
  AOI22D0 U177 ( .A1(\input_value_loc[4][9] ), .A2(n18), .B1(
        \input_value_loc[6][9] ), .B2(n3), .ZN(n148) );
  NR3D0 U178 ( .A1(n8), .A2(n10), .A3(n4), .ZN(n3) );
  NR3D0 U179 ( .A1(n10), .A2(cur_state[1]), .A3(n4), .ZN(n18) );
  AOI22D0 U180 ( .A1(\input_value_loc[2][9] ), .A2(n19), .B1(
        \input_value_loc[3][9] ), .B2(n20), .ZN(n147) );
  NR3D0 U181 ( .A1(n10), .A2(cur_state[2]), .A3(n8), .ZN(n19) );
  AOI22D0 U182 ( .A1(\input_value_loc[0][9] ), .A2(n21), .B1(
        \input_value_loc[1][9] ), .B2(n22), .ZN(n146) );
  CKND0 U183 ( .I(n11), .ZN(n22) );
  CKND2D0 U184 ( .A1(n150), .A2(n4), .ZN(n11) );
  CKND0 U185 ( .I(cur_state[2]), .ZN(n4) );
  NR3D0 U186 ( .A1(cur_state[0]), .A2(cur_state[3]), .A3(n8), .ZN(n150) );
  CKND0 U187 ( .I(cur_state[1]), .ZN(n8) );
  CKND2D0 U188 ( .A1(cur_state[0]), .A2(n9), .ZN(n10) );
  CKND0 U189 ( .I(cur_state[3]), .ZN(n9) );
  NR2D0 U190 ( .A1(cur_state[1]), .A2(cur_state[2]), .ZN(n57) );
endmodule


module routing_engine ( port_dest, control, done );
  input [31:0] port_dest;
  output [19:0] control;
  output done;
  wire   \dst[0][1] , \dst[0][0] , \dst[2][2] , \dst[2][1] , \dst[2][0] ,
         \dst[3][2] , \dst[3][0] , \dst[4][2] , \dst[4][1] , \dst[4][0] ,
         \dst[5][2] , \dst[5][1] , \dst[5][0] , \dst[6][2] , \dst[6][1] ,
         \dst[6][0] , \dst[7][1] , \dst[7][0] , N694, N695, N696, N697, N808,
         N810, N811, N922, N923, N924, N925, N1021, N1022, N1023, N1134, N1135,
         N1136, N1137, N1248, N1249, N1250, N1251, N1362, N1363, N1364, N1365,
         N1446, N1447, N1448, \control[19] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375;
  tri   [19:0] control;
  tri   \control[16] ;
  tri   \control[12] ;
  tri   \control[14] ;
  tri   \control[17] ;
  tri   \control[10] ;
  tri   \control[18] ;
  assign control[13] = \control[19] ;
  assign control[15] = \control[19] ;
  assign control[19] = \control[19] ;

  LHQD1 \dst_reg[0][1]  ( .E(N694), .D(N696), .Q(\dst[0][1] ) );
  LHQD1 \dst_reg[0][0]  ( .E(N694), .D(N695), .Q(\dst[0][0] ) );
  LHD1 \dst_reg[1][1]  ( .E(N808), .D(N810), .QN(n375) );
  LHQD1 \dst_reg[2][2]  ( .E(N922), .D(N925), .Q(\dst[2][2] ) );
  LHQD1 \dst_reg[2][1]  ( .E(N922), .D(N924), .Q(\dst[2][1] ) );
  LHQD1 \dst_reg[2][0]  ( .E(N922), .D(N923), .Q(\dst[2][0] ) );
  LHQD1 \dst_reg[3][2]  ( .E(N1021), .D(N1023), .Q(\dst[3][2] ) );
  LHQD1 \dst_reg[3][0]  ( .E(N1021), .D(N1022), .Q(\dst[3][0] ) );
  LHQD1 \dst_reg[4][2]  ( .E(N1134), .D(N1137), .Q(\dst[4][2] ) );
  LHQD1 \dst_reg[4][1]  ( .E(N1134), .D(N1136), .Q(\dst[4][1] ) );
  LHQD1 \dst_reg[4][0]  ( .E(N1134), .D(N1135), .Q(\dst[4][0] ) );
  LHQD1 \dst_reg[5][2]  ( .E(N1248), .D(N1251), .Q(\dst[5][2] ) );
  LHQD1 \dst_reg[5][1]  ( .E(N1248), .D(N1250), .Q(\dst[5][1] ) );
  LHQD1 \dst_reg[5][0]  ( .E(N1248), .D(N1249), .Q(\dst[5][0] ) );
  LHQD1 \dst_reg[6][2]  ( .E(N1362), .D(N1365), .Q(\dst[6][2] ) );
  LHQD1 \dst_reg[6][1]  ( .E(N1362), .D(N1364), .Q(\dst[6][1] ) );
  LHQD1 \dst_reg[6][0]  ( .E(N1362), .D(N1363), .Q(\dst[6][0] ) );
  LHQD1 \dst_reg[7][1]  ( .E(N1446), .D(N1448), .Q(\dst[7][1] ) );
  LHQD1 \dst_reg[7][0]  ( .E(N1446), .D(N1447), .Q(\dst[7][0] ) );
  LHQD1 \dst_reg[1][2]  ( .E(N808), .D(N811), .Q(control[9]) );
  LHQD1 \dst_reg[0][2]  ( .E(N694), .D(N697), .Q(control[11]) );
  TIEL U448 ( .ZN(\control[19] ) );
  TIEH U449 ( .Z(done) );
  MUX2D0 U450 ( .I0(\dst[2][2] ), .I1(\dst[3][2] ), .S(n1), .Z(control[8]) );
  MUX2ND0 U451 ( .I0(n375), .I1(n2), .S(control[9]), .ZN(control[5]) );
  CKND0 U452 ( .I(n3), .ZN(control[12]) );
  MUX2ND0 U453 ( .I0(n2), .I1(n375), .S(control[9]), .ZN(control[4]) );
  OAI22D0 U454 ( .A1(control[12]), .A2(n4), .B1(n3), .B2(n5), .ZN(n2) );
  MUX2D0 U455 ( .I0(\dst[7][1] ), .I1(\dst[6][1] ), .S(control[16]), .Z(n5) );
  XNR2D0 U456 ( .A1(n6), .A2(control[9]), .ZN(n3) );
  AOI22D0 U457 ( .A1(\dst[5][2] ), .A2(n7), .B1(control[17]), .B2(\dst[4][2] ), 
        .ZN(n6) );
  OA22D0 U458 ( .A1(n7), .A2(\dst[4][1] ), .B1(\dst[5][1] ), .B2(control[17]), 
        .Z(n4) );
  MUX2ND0 U459 ( .I0(n8), .I1(n9), .S(control[7]), .ZN(control[3]) );
  OAI21D0 U460 ( .A1(n10), .A2(n11), .B(n12), .ZN(control[7]) );
  MUX2ND0 U461 ( .I0(n9), .I1(n8), .S(control[7]), .ZN(control[2]) );
  MUX2ND0 U462 ( .I0(\dst[0][0] ), .I1(n13), .S(control[11]), .ZN(n8) );
  OAI22D0 U463 ( .A1(n14), .A2(n15), .B1(control[10]), .B2(n16), .ZN(n9) );
  MUX2ND0 U464 ( .I0(n17), .I1(n18), .S(control[6]), .ZN(control[1]) );
  CKND0 U465 ( .I(n1), .ZN(control[18]) );
  CKND0 U466 ( .I(n15), .ZN(control[10]) );
  CKND0 U467 ( .I(n19), .ZN(control[14]) );
  MUX2ND0 U468 ( .I0(n20), .I1(n21), .S(\dst[6][2] ), .ZN(control[16]) );
  AOI21D0 U469 ( .A1(n22), .A2(\dst[4][2] ), .B(n23), .ZN(n21) );
  MUX2ND0 U470 ( .I0(n24), .I1(n25), .S(\dst[6][1] ), .ZN(n23) );
  AOI21D0 U471 ( .A1(n22), .A2(n26), .B(n27), .ZN(n20) );
  MUX2ND0 U472 ( .I0(n28), .I1(n29), .S(\dst[6][1] ), .ZN(n27) );
  CKND0 U473 ( .I(\dst[4][2] ), .ZN(n26) );
  XNR2D0 U474 ( .A1(\dst[6][1] ), .A2(\dst[4][1] ), .ZN(n22) );
  MUX2ND0 U475 ( .I0(n10), .I1(n30), .S(control[11]), .ZN(control[6]) );
  OA22D0 U476 ( .A1(control[14]), .A2(n31), .B1(n19), .B2(n32), .Z(n10) );
  MUX2ND0 U477 ( .I0(\dst[6][1] ), .I1(\dst[7][1] ), .S(control[16]), .ZN(n32)
         );
  AOI22D0 U478 ( .A1(\dst[4][1] ), .A2(n7), .B1(\dst[5][1] ), .B2(control[17]), 
        .ZN(n31) );
  MUX2ND0 U479 ( .I0(n18), .I1(n17), .S(control[6]), .ZN(control[0]) );
  MUX2ND0 U480 ( .I0(n13), .I1(\dst[0][0] ), .S(control[11]), .ZN(n17) );
  OAI22D0 U481 ( .A1(n33), .A2(control[14]), .B1(n19), .B2(n34), .ZN(n13) );
  MUX2ND0 U482 ( .I0(\dst[6][0] ), .I1(\dst[7][0] ), .S(control[16]), .ZN(n34)
         );
  AOI22D0 U483 ( .A1(\dst[4][0] ), .A2(n7), .B1(\dst[5][0] ), .B2(control[17]), 
        .ZN(n33) );
  OAI22D0 U484 ( .A1(control[10]), .A2(n14), .B1(n16), .B2(n15), .ZN(n18) );
  AOI22D0 U485 ( .A1(\dst[3][2] ), .A2(control[18]), .B1(n1), .B2(\dst[2][2] ), 
        .ZN(n15) );
  OA22D0 U486 ( .A1(\dst[2][0] ), .A2(control[18]), .B1(\dst[3][0] ), .B2(n1), 
        .Z(n16) );
  CKND2D0 U487 ( .A1(n35), .A2(n36), .ZN(n1) );
  CKXOR2D0 U488 ( .A1(control[11]), .A2(n37), .Z(n36) );
  CKXOR2D0 U489 ( .A1(\dst[0][1] ), .A2(n38), .Z(n35) );
  OA22D0 U490 ( .A1(n39), .A2(n19), .B1(control[14]), .B2(n40), .Z(n14) );
  MUX2D0 U491 ( .I0(\dst[6][0] ), .I1(\dst[7][0] ), .S(control[16]), .Z(n40)
         );
  CKXOR2D0 U492 ( .A1(n41), .A2(n11), .Z(n19) );
  AOI22D0 U493 ( .A1(\dst[4][2] ), .A2(n7), .B1(control[17]), .B2(\dst[5][2] ), 
        .ZN(n41) );
  OA22D0 U494 ( .A1(n7), .A2(\dst[5][0] ), .B1(control[17]), .B2(\dst[4][0] ), 
        .Z(n39) );
  CKND0 U495 ( .I(control[17]), .ZN(n7) );
  MUX4ND0 U496 ( .I0(n28), .I1(n29), .I2(n24), .I3(n25), .S0(\dst[4][1] ), 
        .S1(\dst[4][2] ), .ZN(control[17]) );
  AOI22D0 U497 ( .A1(\dst[2][2] ), .A2(\dst[2][1] ), .B1(control[11]), .B2(
        \dst[0][1] ), .ZN(n25) );
  AOI22D0 U498 ( .A1(n38), .A2(\dst[2][2] ), .B1(n30), .B2(control[11]), .ZN(
        n24) );
  OA21D0 U499 ( .A1(\dst[2][2] ), .A2(n38), .B(n12), .Z(n29) );
  CKND2D0 U500 ( .A1(\dst[0][1] ), .A2(n11), .ZN(n12) );
  AOI22D0 U501 ( .A1(n38), .A2(n37), .B1(n11), .B2(n30), .ZN(n28) );
  CKND0 U502 ( .I(\dst[0][1] ), .ZN(n30) );
  CKND0 U503 ( .I(control[11]), .ZN(n11) );
  CKND0 U504 ( .I(\dst[2][2] ), .ZN(n37) );
  CKND0 U505 ( .I(\dst[2][1] ), .ZN(n38) );
  OAI211D0 U506 ( .A1(port_dest[23]), .A2(n42), .B(n43), .C(n44), .ZN(N925) );
  AOI21D0 U507 ( .A1(n45), .A2(port_dest[22]), .B(n46), .ZN(n42) );
  OAI221D0 U508 ( .A1(n47), .A2(n48), .B1(port_dest[23]), .B2(n49), .C(n44), 
        .ZN(N924) );
  AOI21D0 U509 ( .A1(n50), .A2(n51), .B(n52), .ZN(n44) );
  CKND0 U510 ( .I(n53), .ZN(n52) );
  NR2D0 U511 ( .A1(n54), .A2(n55), .ZN(n49) );
  AOI21D0 U512 ( .A1(n56), .A2(n57), .B(port_dest[23]), .ZN(n47) );
  CKND2D0 U513 ( .A1(n58), .A2(n53), .ZN(N923) );
  ND3D0 U514 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n53) );
  MUX2ND0 U515 ( .I0(n62), .I1(port_dest[20]), .S(port_dest[23]), .ZN(n58) );
  AOI21D0 U516 ( .A1(n63), .A2(n64), .B(n51), .ZN(n62) );
  OAI21D0 U517 ( .A1(n65), .A2(n54), .B(n66), .ZN(n64) );
  INR3D0 U518 ( .A1(n67), .B1(n68), .B2(n69), .ZN(n54) );
  AOI211D0 U519 ( .A1(n70), .A2(n71), .B(n72), .C(n55), .ZN(n65) );
  ND4D0 U520 ( .A1(n57), .A2(n69), .A3(n56), .A4(n73), .ZN(N922) );
  NR4D0 U521 ( .A1(port_dest[23]), .A2(n55), .A3(n51), .A4(n59), .ZN(n73) );
  CKND0 U522 ( .I(n74), .ZN(n59) );
  NR3D0 U523 ( .A1(n60), .A2(n75), .A3(n76), .ZN(n51) );
  NR2D0 U524 ( .A1(n67), .A2(n68), .ZN(n55) );
  CKND0 U525 ( .I(n57), .ZN(n68) );
  CKND0 U526 ( .I(n46), .ZN(n56) );
  CKND2D0 U527 ( .A1(n63), .A2(n66), .ZN(n46) );
  CKND2D0 U528 ( .A1(n77), .A2(n45), .ZN(n66) );
  CKND0 U529 ( .I(n78), .ZN(n45) );
  CKND2D0 U530 ( .A1(n75), .A2(n79), .ZN(n63) );
  OAI21D0 U531 ( .A1(port_dest[27]), .A2(n80), .B(n81), .ZN(N811) );
  AOI221D0 U532 ( .A1(n82), .A2(n83), .B1(n84), .B2(port_dest[26]), .C(n85), 
        .ZN(n80) );
  OAI222D0 U533 ( .A1(n86), .A2(n87), .B1(n88), .B2(n89), .C1(n90), .C2(n91), 
        .ZN(N810) );
  NR2D0 U534 ( .A1(n82), .A2(n92), .ZN(n88) );
  AOI21D0 U535 ( .A1(n93), .A2(n94), .B(port_dest[27]), .ZN(n86) );
  IND3D0 U536 ( .A1(n85), .B1(n95), .B2(n96), .ZN(N808) );
  CKND0 U537 ( .I(n82), .ZN(n96) );
  IOA21D0 U538 ( .A1(n83), .A2(n92), .B(n93), .ZN(n85) );
  AOI22D0 U539 ( .A1(n84), .A2(n97), .B1(n83), .B2(n98), .ZN(n93) );
  CKND0 U540 ( .I(n99), .ZN(n84) );
  OAI211D0 U541 ( .A1(port_dest[31]), .A2(n100), .B(n101), .C(n102), .ZN(N697)
         );
  AOI211D0 U542 ( .A1(n103), .A2(port_dest[30]), .B(n104), .C(n105), .ZN(n100)
         );
  OAI221D0 U543 ( .A1(n106), .A2(n107), .B1(port_dest[31]), .B2(n108), .C(n101), .ZN(N696) );
  OA31D0 U544 ( .A1(n109), .A2(n110), .A3(n104), .B(n111), .Z(n106) );
  CKND2D0 U545 ( .A1(n112), .A2(n101), .ZN(N695) );
  IND2D0 U546 ( .A1(n113), .B1(n114), .ZN(n101) );
  MUX2ND0 U547 ( .I0(n115), .I1(port_dest[28]), .S(port_dest[31]), .ZN(n112)
         );
  NR2D0 U548 ( .A1(n105), .A2(n116), .ZN(n115) );
  MAOI22D0 U549 ( .A1(n117), .A2(n118), .B1(n119), .B2(n120), .ZN(n116) );
  OAI32D0 U550 ( .A1(n121), .A2(n122), .A3(n109), .B1(n123), .B2(n124), .ZN(
        n117) );
  NR2D0 U551 ( .A1(n110), .A2(port_dest[28]), .ZN(n121) );
  ND4D0 U552 ( .A1(n113), .A2(n125), .A3(n126), .A4(n127), .ZN(N694) );
  INR2D0 U553 ( .A1(n108), .B1(n104), .ZN(n127) );
  OAI21D0 U554 ( .A1(n120), .A2(n119), .B(n118), .ZN(n104) );
  IND2D0 U555 ( .A1(n128), .B1(n103), .ZN(n118) );
  AOI211D0 U556 ( .A1(n129), .A2(n130), .B(n122), .C(n105), .ZN(n108) );
  INR3D0 U557 ( .A1(n119), .B1(n120), .B2(n131), .ZN(n105) );
  NR3D0 U558 ( .A1(n109), .A2(n110), .A3(n132), .ZN(n122) );
  CKND0 U559 ( .I(n125), .ZN(n110) );
  CKND2D0 U560 ( .A1(n133), .A2(n134), .ZN(N1448) );
  OAI31D0 U561 ( .A1(n135), .A2(n136), .A3(n137), .B(n138), .ZN(n134) );
  CKND0 U562 ( .I(n139), .ZN(n137) );
  AOI211D0 U563 ( .A1(n140), .A2(n141), .B(n142), .C(n143), .ZN(n135) );
  CKND0 U564 ( .I(n144), .ZN(n143) );
  CKND2D0 U565 ( .A1(n145), .A2(port_dest[1]), .ZN(n141) );
  MUX2ND0 U566 ( .I0(n146), .I1(n147), .S(port_dest[3]), .ZN(N1447) );
  AOI21D0 U567 ( .A1(n148), .A2(n139), .B(n136), .ZN(n146) );
  ND3D0 U568 ( .A1(n149), .A2(n150), .A3(n151), .ZN(n139) );
  OAI21D0 U569 ( .A1(n142), .A2(n152), .B(n144), .ZN(n148) );
  CKND2D0 U570 ( .A1(n153), .A2(n149), .ZN(n144) );
  AOI32D0 U571 ( .A1(n154), .A2(n155), .A3(n156), .B1(n157), .B2(n158), .ZN(
        n152) );
  OAI21D0 U572 ( .A1(n159), .A2(n160), .B(n147), .ZN(n156) );
  ND4D0 U573 ( .A1(n145), .A2(n150), .A3(n140), .A4(n161), .ZN(N1446) );
  NR4D0 U574 ( .A1(port_dest[3]), .A2(n142), .A3(n136), .A4(n151), .ZN(n161)
         );
  IINR4D0 U575 ( .A1(n162), .A2(n163), .B1(n151), .B2(n153), .ZN(n136) );
  AOI21D0 U576 ( .A1(n164), .A2(n165), .B(n166), .ZN(n151) );
  INR2D0 U577 ( .A1(n149), .B1(n167), .ZN(n162) );
  AOI211D0 U578 ( .A1(n168), .A2(n169), .B(n157), .C(n170), .ZN(n149) );
  CKND0 U579 ( .I(n171), .ZN(n157) );
  AN4D0 U580 ( .A1(n158), .A2(n169), .A3(n171), .A4(n168), .Z(n142) );
  CKND0 U581 ( .I(n170), .ZN(n158) );
  OA21D0 U582 ( .A1(n170), .A2(n171), .B(n154), .Z(n140) );
  ND3D0 U583 ( .A1(n172), .A2(n173), .A3(n145), .ZN(n154) );
  OAI21D0 U584 ( .A1(port_dest[7]), .A2(n174), .B(n175), .ZN(n171) );
  OAI21D0 U585 ( .A1(n176), .A2(n177), .B(n145), .ZN(n170) );
  CKND0 U586 ( .I(n153), .ZN(n150) );
  NR2D0 U587 ( .A1(n164), .A2(n165), .ZN(n153) );
  OA21D0 U588 ( .A1(n159), .A2(n160), .B(n155), .Z(n145) );
  CKND2D0 U589 ( .A1(n178), .A2(port_dest[7]), .ZN(n155) );
  OAI221D0 U590 ( .A1(port_dest[7]), .A2(n179), .B1(n180), .B2(n168), .C(n181), 
        .ZN(N1365) );
  NR2D0 U591 ( .A1(n182), .A2(n183), .ZN(n181) );
  ND3D0 U592 ( .A1(n184), .A2(n185), .A3(n186), .ZN(n168) );
  NR2D0 U593 ( .A1(n187), .A2(n188), .ZN(n179) );
  OAI221D0 U594 ( .A1(n189), .A2(n190), .B1(port_dest[7]), .B2(n191), .C(n192), 
        .ZN(N1364) );
  AOI21D0 U595 ( .A1(n193), .A2(n194), .B(port_dest[7]), .ZN(n189) );
  CKND2D0 U596 ( .A1(n195), .A2(n192), .ZN(N1363) );
  CKND0 U597 ( .I(n183), .ZN(n192) );
  NR2D0 U598 ( .A1(n163), .A2(n167), .ZN(n183) );
  ND3D0 U599 ( .A1(n164), .A2(n166), .A3(n165), .ZN(n163) );
  NR2D0 U600 ( .A1(n196), .A2(port_dest[7]), .ZN(n165) );
  MUX2ND0 U601 ( .I0(n197), .I1(port_dest[4]), .S(port_dest[7]), .ZN(n195) );
  NR2D0 U602 ( .A1(n187), .A2(n198), .ZN(n197) );
  AOI22D0 U603 ( .A1(n199), .A2(n200), .B1(n201), .B2(n202), .ZN(n198) );
  OAI32D0 U604 ( .A1(n203), .A2(n178), .A3(n204), .B1(n174), .B2(n184), .ZN(
        n199) );
  NR2D0 U605 ( .A1(n205), .A2(port_dest[4]), .ZN(n203) );
  ND4D0 U606 ( .A1(n176), .A2(n191), .A3(n193), .A4(n167), .ZN(N1362) );
  IND2D0 U607 ( .A1(n206), .B1(n207), .ZN(n167) );
  CKND0 U608 ( .I(n188), .ZN(n193) );
  OAI21D0 U609 ( .A1(n196), .A2(n164), .B(n200), .ZN(n188) );
  ND3D0 U610 ( .A1(n186), .A2(n184), .A3(n169), .ZN(n200) );
  CKND0 U611 ( .I(n175), .ZN(n184) );
  CKND0 U612 ( .I(n201), .ZN(n164) );
  AOI211D0 U613 ( .A1(n186), .A2(n175), .B(n187), .C(n204), .ZN(n191) );
  AN2D0 U614 ( .A1(n194), .A2(n172), .Z(n204) );
  NR3D0 U615 ( .A1(n196), .A2(n201), .A3(n166), .ZN(n187) );
  CKND2D0 U616 ( .A1(n208), .A2(n209), .ZN(n166) );
  AOI21D0 U617 ( .A1(n210), .A2(n211), .B(n212), .ZN(n201) );
  CKND0 U618 ( .I(n202), .ZN(n196) );
  NR3D0 U619 ( .A1(n175), .A2(n169), .A3(n174), .ZN(n202) );
  NR2D0 U620 ( .A1(n210), .A2(n211), .ZN(n169) );
  AOI21D0 U621 ( .A1(n213), .A2(n214), .B(n215), .ZN(n175) );
  CKND0 U622 ( .I(n174), .ZN(n186) );
  CKND2D0 U623 ( .A1(n194), .A2(n177), .ZN(n174) );
  CKND0 U624 ( .I(n172), .ZN(n177) );
  NR2D0 U625 ( .A1(n216), .A2(n217), .ZN(n172) );
  NR2D0 U626 ( .A1(n178), .A2(n205), .ZN(n194) );
  CKND0 U627 ( .I(n173), .ZN(n176) );
  CKND2D0 U628 ( .A1(n159), .A2(n160), .ZN(n173) );
  CKND0 U629 ( .I(n205), .ZN(n160) );
  AOI21D0 U630 ( .A1(n218), .A2(n213), .B(n219), .ZN(n205) );
  NR2D0 U631 ( .A1(port_dest[7]), .A2(n178), .ZN(n159) );
  NR2D0 U632 ( .A1(n218), .A2(n213), .ZN(n178) );
  OAI221D0 U633 ( .A1(n220), .A2(n221), .B1(port_dest[11]), .B2(n222), .C(n223), .ZN(N1251) );
  NR2D0 U634 ( .A1(n224), .A2(port_dest[11]), .ZN(n220) );
  OAI211D0 U635 ( .A1(port_dest[11]), .A2(n225), .B(n226), .C(n223), .ZN(N1250) );
  AOI21D0 U636 ( .A1(n227), .A2(n228), .B(n229), .ZN(n225) );
  OAI21D0 U637 ( .A1(n230), .A2(n231), .B(n232), .ZN(n228) );
  CKND0 U638 ( .I(port_dest[9]), .ZN(n230) );
  CKND2D0 U639 ( .A1(n233), .A2(n223), .ZN(N1249) );
  CKND2D0 U640 ( .A1(n206), .A2(n207), .ZN(n223) );
  NR2D0 U641 ( .A1(n209), .A2(n208), .ZN(n206) );
  ND3D0 U642 ( .A1(n210), .A2(n212), .A3(n211), .ZN(n209) );
  NR2D0 U643 ( .A1(n234), .A2(port_dest[11]), .ZN(n211) );
  MUX2ND0 U644 ( .I0(n235), .I1(port_dest[8]), .S(port_dest[11]), .ZN(n233) );
  AOI21D0 U645 ( .A1(n236), .A2(n237), .B(n229), .ZN(n235) );
  OAI22D0 U646 ( .A1(n234), .A2(n210), .B1(n238), .B2(n239), .ZN(n236) );
  AOI211D0 U647 ( .A1(n219), .A2(n240), .B(n241), .C(n242), .ZN(n239) );
  CKND0 U648 ( .I(n218), .ZN(n241) );
  IND4D0 U649 ( .A1(n207), .B1(n217), .B2(n222), .B3(n232), .ZN(N1248) );
  NR2D0 U650 ( .A1(n238), .A2(n242), .ZN(n232) );
  NR2D0 U651 ( .A1(n216), .A2(n231), .ZN(n242) );
  CKND0 U652 ( .I(n243), .ZN(n216) );
  INR2D0 U653 ( .A1(n214), .B1(n215), .ZN(n238) );
  INR2D0 U654 ( .A1(n227), .B1(n229), .ZN(n222) );
  AN4D0 U655 ( .A1(n208), .A2(n224), .A3(n210), .A4(n212), .Z(n229) );
  CKND0 U656 ( .I(n244), .ZN(n212) );
  AOI21D0 U657 ( .A1(n245), .A2(n246), .B(n247), .ZN(n208) );
  OA21D0 U658 ( .A1(n234), .A2(n210), .B(n237), .Z(n227) );
  ND3D0 U659 ( .A1(n224), .A2(n210), .A3(n244), .ZN(n237) );
  NR2D0 U660 ( .A1(n245), .A2(n246), .ZN(n244) );
  CKND0 U661 ( .I(n234), .ZN(n224) );
  OAI21D0 U662 ( .A1(port_dest[15]), .A2(n248), .B(n249), .ZN(n210) );
  CKND2D0 U663 ( .A1(n214), .A2(n215), .ZN(n234) );
  AO21D0 U664 ( .A1(n250), .A2(n251), .B(n252), .Z(n215) );
  NR2D0 U665 ( .A1(n231), .A2(n243), .ZN(n214) );
  NR2D0 U666 ( .A1(n253), .A2(n254), .ZN(n243) );
  NR2D0 U667 ( .A1(n231), .A2(port_dest[11]), .ZN(n217) );
  CKND2D0 U668 ( .A1(n218), .A2(n219), .ZN(n231) );
  OAI21D0 U669 ( .A1(port_dest[15]), .A2(n255), .B(n256), .ZN(n219) );
  CKND2D0 U670 ( .A1(n255), .A2(port_dest[15]), .ZN(n218) );
  NR2D0 U671 ( .A1(n257), .A2(n258), .ZN(n207) );
  OAI211D0 U672 ( .A1(port_dest[15]), .A2(n259), .B(n260), .C(n261), .ZN(N1137) );
  CKND0 U673 ( .I(n262), .ZN(n261) );
  OA21D0 U674 ( .A1(n248), .A2(n263), .B(n264), .Z(n259) );
  OAI221D0 U675 ( .A1(port_dest[15]), .A2(n265), .B1(n266), .B2(n267), .C(n260), .ZN(N1136) );
  MOAI22D0 U676 ( .A1(port_dest[15]), .A2(n268), .B1(n246), .B2(n269), .ZN(
        n267) );
  NR2D0 U677 ( .A1(n270), .A2(n271), .ZN(n268) );
  INR2D0 U678 ( .A1(n272), .B1(n273), .ZN(n265) );
  OAI221D0 U679 ( .A1(n273), .A2(n274), .B1(n250), .B2(n275), .C(n260), .ZN(
        N1135) );
  IND2D0 U680 ( .A1(n257), .B1(n258), .ZN(n260) );
  AN3D0 U681 ( .A1(n247), .A2(n245), .A3(n246), .Z(n258) );
  AOI32D0 U682 ( .A1(n276), .A2(n250), .A3(n277), .B1(n269), .B2(n246), .ZN(
        n274) );
  NR2D0 U683 ( .A1(n278), .A2(port_dest[15]), .ZN(n246) );
  OAI32D0 U684 ( .A1(n279), .A2(n255), .A3(n280), .B1(n281), .B2(n252), .ZN(
        n277) );
  CKND0 U685 ( .I(n282), .ZN(n255) );
  NR2D0 U686 ( .A1(n256), .A2(port_dest[12]), .ZN(n279) );
  CKND0 U687 ( .I(n270), .ZN(n276) );
  ND4D0 U688 ( .A1(n254), .A2(n272), .A3(n264), .A4(n257), .ZN(N1134) );
  OAI31D0 U689 ( .A1(n283), .A2(port_dest[19]), .A3(n284), .B(n285), .ZN(n257)
         );
  AOI211D0 U690 ( .A1(n286), .A2(n269), .B(n270), .C(n273), .ZN(n264) );
  NR3D0 U691 ( .A1(n278), .A2(n269), .A3(n247), .ZN(n273) );
  OAI21D0 U692 ( .A1(port_dest[19]), .A2(n283), .B(n284), .ZN(n247) );
  CKND0 U693 ( .I(n286), .ZN(n278) );
  NR2D0 U694 ( .A1(n287), .A2(n248), .ZN(n270) );
  CKND0 U695 ( .I(n245), .ZN(n269) );
  OAI21D0 U696 ( .A1(n288), .A2(n289), .B(n290), .ZN(n245) );
  NR2D0 U697 ( .A1(n248), .A2(n249), .ZN(n286) );
  CKND0 U698 ( .I(n287), .ZN(n249) );
  CKND2D0 U699 ( .A1(n288), .A2(n289), .ZN(n287) );
  CKND2D0 U700 ( .A1(n251), .A2(n252), .ZN(n248) );
  IAO21D0 U701 ( .A1(n281), .A2(n252), .B(n280), .ZN(n272) );
  NR2D0 U702 ( .A1(n253), .A2(n271), .ZN(n280) );
  OAI21D0 U703 ( .A1(n291), .A2(n292), .B(n293), .ZN(n252) );
  CKND0 U704 ( .I(n251), .ZN(n281) );
  INR2D0 U705 ( .A1(n253), .B1(n271), .ZN(n251) );
  CKND2D0 U706 ( .A1(n291), .A2(n292), .ZN(n253) );
  ND3D0 U707 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n292) );
  NR2D0 U708 ( .A1(n271), .A2(port_dest[15]), .ZN(n254) );
  IND2D0 U709 ( .A1(n256), .B1(n282), .ZN(n271) );
  CKND2D0 U710 ( .A1(n297), .A2(port_dest[19]), .ZN(n282) );
  AOI21D0 U711 ( .A1(n294), .A2(n295), .B(n296), .ZN(n256) );
  OAI221D0 U712 ( .A1(n298), .A2(n289), .B1(port_dest[19]), .B2(n299), .C(n300), .ZN(N1023) );
  CKND0 U713 ( .I(port_dest[18]), .ZN(n298) );
  MUX2ND0 U714 ( .I0(n301), .I1(n302), .S(port_dest[19]), .ZN(N1022) );
  INR2D0 U715 ( .A1(n303), .B1(n304), .ZN(n301) );
  AOI21D0 U716 ( .A1(n284), .A2(n305), .B(n306), .ZN(n304) );
  AOI31D0 U717 ( .A1(n307), .A2(n308), .A3(n290), .B(n309), .ZN(n306) );
  AOI221D0 U718 ( .A1(n288), .A2(n307), .B1(n310), .B2(n296), .C(n297), .ZN(
        n309) );
  OAI21D0 U719 ( .A1(port_dest[16]), .A2(n293), .B(n311), .ZN(n310) );
  CKND0 U720 ( .I(n291), .ZN(n311) );
  IND2D0 U721 ( .A1(n289), .B1(n299), .ZN(N1021) );
  AN2D0 U722 ( .A1(n303), .A2(n312), .Z(n299) );
  OAI31D0 U723 ( .A1(n288), .A2(n284), .A3(n290), .B(n307), .ZN(n312) );
  CKND0 U724 ( .I(n313), .ZN(n290) );
  CKND0 U725 ( .I(n308), .ZN(n288) );
  IND3D0 U726 ( .A1(n284), .B1(n305), .B2(n285), .ZN(n303) );
  AOI21D0 U727 ( .A1(n60), .A2(n61), .B(n74), .ZN(n285) );
  OAI21D0 U728 ( .A1(n92), .A2(n89), .B(n82), .ZN(n74) );
  NR2D0 U729 ( .A1(n113), .A2(n114), .ZN(n82) );
  INR2D0 U730 ( .A1(n131), .B1(n314), .ZN(n114) );
  ND4D0 U731 ( .A1(n315), .A2(n316), .A3(n317), .A4(n318), .ZN(n113) );
  AOI33D0 U732 ( .A1(n319), .A2(port_dest[10]), .A3(port_dest[8]), .B1(n320), 
        .B2(port_dest[2]), .B3(port_dest[0]), .ZN(n318) );
  AOI33D0 U733 ( .A1(port_dest[12]), .A2(n262), .A3(port_dest[13]), .B1(
        port_dest[16]), .B2(n321), .B3(port_dest[17]), .ZN(n317) );
  AOI33D0 U734 ( .A1(port_dest[4]), .A2(n182), .A3(port_dest[5]), .B1(
        port_dest[28]), .B2(n322), .B3(port_dest[29]), .ZN(n316) );
  AOI33D0 U735 ( .A1(port_dest[20]), .A2(n323), .A3(port_dest[21]), .B1(
        port_dest[24]), .B2(n324), .B3(port_dest[25]), .ZN(n315) );
  CKND0 U736 ( .I(n283), .ZN(n305) );
  ND3D0 U737 ( .A1(n308), .A2(n313), .A3(n307), .ZN(n283) );
  OAI21D0 U738 ( .A1(port_dest[23]), .A2(n76), .B(n75), .ZN(n313) );
  OAI21D0 U739 ( .A1(port_dest[23]), .A2(n78), .B(n77), .ZN(n308) );
  NR2D0 U740 ( .A1(n60), .A2(n61), .ZN(n284) );
  NR3D0 U741 ( .A1(n75), .A2(port_dest[23]), .A3(n76), .ZN(n61) );
  CKND0 U742 ( .I(n79), .ZN(n76) );
  NR2D0 U743 ( .A1(n78), .A2(n77), .ZN(n79) );
  INR2D0 U744 ( .A1(n97), .B1(n95), .ZN(n77) );
  NR2D0 U745 ( .A1(n99), .A2(port_dest[27]), .ZN(n95) );
  ND3D0 U746 ( .A1(n69), .A2(n67), .A3(n57), .ZN(n78) );
  AOI21D0 U747 ( .A1(n325), .A2(n83), .B(n326), .ZN(n75) );
  CKND2D0 U748 ( .A1(n92), .A2(n89), .ZN(n60) );
  ND3D0 U749 ( .A1(n326), .A2(n325), .A3(n83), .ZN(n89) );
  NR2D0 U750 ( .A1(n99), .A2(n97), .ZN(n83) );
  AOI21D0 U751 ( .A1(n111), .A2(n103), .B(n128), .ZN(n97) );
  CKND2D0 U752 ( .A1(n94), .A2(n90), .ZN(n99) );
  NR2D0 U753 ( .A1(n327), .A2(n328), .ZN(n90) );
  CKND0 U754 ( .I(n98), .ZN(n326) );
  NR2D0 U755 ( .A1(n119), .A2(n329), .ZN(n98) );
  INR2D0 U756 ( .A1(n314), .B1(n131), .ZN(n92) );
  ND4D0 U757 ( .A1(n330), .A2(n331), .A3(n332), .A4(n333), .ZN(n131) );
  AOI33D0 U758 ( .A1(port_dest[10]), .A2(n240), .A3(n319), .B1(port_dest[2]), 
        .B2(n147), .B3(n320), .ZN(n333) );
  AOI33D0 U759 ( .A1(n262), .A2(n275), .A3(port_dest[13]), .B1(n321), .B2(n302), .B3(port_dest[17]), .ZN(n332) );
  AOI33D0 U760 ( .A1(n182), .A2(n334), .A3(port_dest[5]), .B1(n322), .B2(n335), 
        .B3(port_dest[29]), .ZN(n331) );
  AOI33D0 U761 ( .A1(n323), .A2(n70), .A3(port_dest[21]), .B1(n324), .B2(n336), 
        .B3(port_dest[25]), .ZN(n330) );
  CKND2D0 U762 ( .A1(n329), .A2(n119), .ZN(n314) );
  ND4D0 U763 ( .A1(n337), .A2(n338), .A3(n339), .A4(n340), .ZN(n119) );
  AOI33D0 U764 ( .A1(port_dest[10]), .A2(n341), .A3(port_dest[8]), .B1(
        port_dest[2]), .B2(n342), .B3(port_dest[0]), .ZN(n340) );
  AOI33D0 U765 ( .A1(n262), .A2(n266), .A3(port_dest[12]), .B1(n321), .B2(n343), .B3(port_dest[16]), .ZN(n339) );
  AOI33D0 U766 ( .A1(n182), .A2(n190), .A3(port_dest[4]), .B1(n322), .B2(n107), 
        .B3(port_dest[28]), .ZN(n338) );
  AOI33D0 U767 ( .A1(n323), .A2(n48), .A3(port_dest[20]), .B1(n324), .B2(n87), 
        .B3(port_dest[24]), .ZN(n337) );
  NR2D0 U768 ( .A1(n120), .A2(port_dest[31]), .ZN(n329) );
  CKND2D0 U769 ( .A1(n103), .A2(n128), .ZN(n120) );
  ND4D0 U770 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .ZN(n128) );
  AOI33D0 U771 ( .A1(n341), .A2(n240), .A3(port_dest[10]), .B1(n342), .B2(n147), .B3(port_dest[2]), .ZN(n347) );
  AOI33D0 U772 ( .A1(n275), .A2(n266), .A3(n262), .B1(n302), .B2(n343), .B3(
        n321), .ZN(n346) );
  CKND0 U773 ( .I(n300), .ZN(n321) );
  CKND2D0 U774 ( .A1(port_dest[19]), .A2(port_dest[18]), .ZN(n300) );
  NR2D0 U775 ( .A1(n250), .A2(n263), .ZN(n262) );
  CKND0 U776 ( .I(port_dest[14]), .ZN(n263) );
  AOI33D0 U777 ( .A1(n334), .A2(n190), .A3(n182), .B1(n335), .B2(n107), .B3(
        n322), .ZN(n345) );
  CKND0 U778 ( .I(n102), .ZN(n322) );
  CKND2D0 U779 ( .A1(port_dest[31]), .A2(port_dest[30]), .ZN(n102) );
  NR2D0 U780 ( .A1(n185), .A2(n180), .ZN(n182) );
  CKND0 U781 ( .I(port_dest[6]), .ZN(n180) );
  AOI33D0 U782 ( .A1(n70), .A2(n48), .A3(n323), .B1(n336), .B2(n87), .B3(n324), 
        .ZN(n344) );
  CKND0 U783 ( .I(n81), .ZN(n324) );
  CKND2D0 U784 ( .A1(port_dest[27]), .A2(port_dest[26]), .ZN(n81) );
  CKND0 U785 ( .I(n43), .ZN(n323) );
  CKND2D0 U786 ( .A1(port_dest[23]), .A2(port_dest[22]), .ZN(n43) );
  NR2D0 U787 ( .A1(n123), .A2(n130), .ZN(n103) );
  CKND0 U788 ( .I(n124), .ZN(n130) );
  CKND2D0 U789 ( .A1(n307), .A2(n295), .ZN(n289) );
  INR4D0 U790 ( .A1(n296), .B1(n293), .B2(n297), .B3(n291), .ZN(n307) );
  AOI21D0 U791 ( .A1(n50), .A2(n57), .B(n67), .ZN(n291) );
  CKND0 U792 ( .I(n294), .ZN(n297) );
  CKND2D0 U793 ( .A1(n72), .A2(port_dest[23]), .ZN(n294) );
  AOI31D0 U794 ( .A1(n57), .A2(n50), .A3(n67), .B(n69), .ZN(n293) );
  OAI21D0 U795 ( .A1(n328), .A2(n91), .B(n327), .ZN(n69) );
  AOI21D0 U796 ( .A1(n111), .A2(n129), .B(n124), .ZN(n327) );
  ND4D0 U797 ( .A1(n348), .A2(n349), .A3(n350), .A4(n351), .ZN(n124) );
  AOI33D0 U798 ( .A1(port_dest[16]), .A2(n352), .A3(port_dest[17]), .B1(
        port_dest[12]), .B2(n353), .B3(port_dest[13]), .ZN(n351) );
  AOI33D0 U799 ( .A1(port_dest[4]), .A2(n354), .A3(port_dest[5]), .B1(
        port_dest[24]), .B2(n355), .B3(port_dest[25]), .ZN(n350) );
  AOI33D0 U800 ( .A1(port_dest[28]), .A2(n356), .A3(port_dest[29]), .B1(
        port_dest[20]), .B2(n357), .B3(port_dest[21]), .ZN(n349) );
  AOI33D0 U801 ( .A1(n319), .A2(n221), .A3(port_dest[8]), .B1(n320), .B2(n358), 
        .B3(port_dest[0]), .ZN(n348) );
  CKND0 U802 ( .I(n123), .ZN(n129) );
  ND3D0 U803 ( .A1(n359), .A2(n125), .A3(n132), .ZN(n123) );
  CKND2D0 U804 ( .A1(n328), .A2(n91), .ZN(n67) );
  CKND2D0 U805 ( .A1(n94), .A2(n325), .ZN(n91) );
  AOI21D0 U806 ( .A1(port_dest[31]), .A2(n109), .B(n360), .ZN(n94) );
  AOI21D0 U807 ( .A1(n125), .A2(n126), .B(n132), .ZN(n328) );
  ND4D0 U808 ( .A1(n361), .A2(n362), .A3(n363), .A4(n364), .ZN(n132) );
  AOI33D0 U809 ( .A1(n352), .A2(n302), .A3(port_dest[17]), .B1(n353), .B2(n275), .B3(port_dest[13]), .ZN(n364) );
  AOI33D0 U810 ( .A1(n354), .A2(n334), .A3(port_dest[5]), .B1(n355), .B2(n336), 
        .B3(port_dest[25]), .ZN(n363) );
  AOI33D0 U811 ( .A1(n356), .A2(n335), .A3(port_dest[29]), .B1(n357), .B2(n70), 
        .B3(port_dest[21]), .ZN(n362) );
  AOI33D0 U812 ( .A1(n221), .A2(n240), .A3(n319), .B1(n147), .B2(n358), .B3(
        n320), .ZN(n361) );
  CKND0 U813 ( .I(n133), .ZN(n320) );
  CKND2D0 U814 ( .A1(port_dest[1]), .A2(port_dest[3]), .ZN(n133) );
  CKND0 U815 ( .I(n226), .ZN(n319) );
  CKND2D0 U816 ( .A1(port_dest[9]), .A2(port_dest[11]), .ZN(n226) );
  NR2D0 U817 ( .A1(n72), .A2(n365), .ZN(n57) );
  OAI21D0 U818 ( .A1(port_dest[23]), .A2(n72), .B(n365), .ZN(n296) );
  CKND0 U819 ( .I(n71), .ZN(n365) );
  OAI21D0 U820 ( .A1(n366), .A2(port_dest[27]), .B(n360), .ZN(n71) );
  NR2D0 U821 ( .A1(n125), .A2(n126), .ZN(n360) );
  NR2D0 U822 ( .A1(port_dest[31]), .A2(n109), .ZN(n126) );
  CKND0 U823 ( .I(n359), .ZN(n109) );
  ND4D0 U824 ( .A1(n367), .A2(n368), .A3(n369), .A4(n370), .ZN(n125) );
  AOI33D0 U825 ( .A1(n352), .A2(n343), .A3(port_dest[16]), .B1(n353), .B2(n266), .B3(port_dest[12]), .ZN(n370) );
  AOI33D0 U826 ( .A1(n341), .A2(n221), .A3(port_dest[8]), .B1(n354), .B2(n190), 
        .B3(port_dest[4]), .ZN(n369) );
  AOI33D0 U827 ( .A1(n342), .A2(n358), .A3(port_dest[0]), .B1(n355), .B2(n87), 
        .B3(port_dest[24]), .ZN(n368) );
  AOI33D0 U828 ( .A1(n356), .A2(n107), .A3(port_dest[28]), .B1(n357), .B2(n48), 
        .B3(port_dest[20]), .ZN(n367) );
  NR2D0 U829 ( .A1(n111), .A2(n359), .ZN(n366) );
  NR3D0 U830 ( .A1(n325), .A2(n111), .A3(n359), .ZN(n72) );
  ND4D0 U831 ( .A1(n371), .A2(n372), .A3(n373), .A4(n374), .ZN(n359) );
  AOI33D0 U832 ( .A1(n302), .A2(n343), .A3(n352), .B1(n275), .B2(n266), .B3(
        n353), .ZN(n374) );
  NR2D0 U833 ( .A1(n250), .A2(port_dest[14]), .ZN(n353) );
  CKND0 U834 ( .I(port_dest[15]), .ZN(n250) );
  CKND0 U835 ( .I(port_dest[13]), .ZN(n266) );
  CKND0 U836 ( .I(port_dest[12]), .ZN(n275) );
  NR2D0 U837 ( .A1(n295), .A2(port_dest[18]), .ZN(n352) );
  CKND0 U838 ( .I(port_dest[19]), .ZN(n295) );
  CKND0 U839 ( .I(port_dest[17]), .ZN(n343) );
  CKND0 U840 ( .I(port_dest[16]), .ZN(n302) );
  AOI33D0 U841 ( .A1(n221), .A2(n240), .A3(n341), .B1(n334), .B2(n190), .B3(
        n354), .ZN(n373) );
  NR2D0 U842 ( .A1(n185), .A2(port_dest[6]), .ZN(n354) );
  CKND0 U843 ( .I(port_dest[7]), .ZN(n185) );
  CKND0 U844 ( .I(port_dest[5]), .ZN(n190) );
  CKND0 U845 ( .I(port_dest[4]), .ZN(n334) );
  NR2D0 U846 ( .A1(n213), .A2(port_dest[9]), .ZN(n341) );
  CKND0 U847 ( .I(port_dest[11]), .ZN(n213) );
  CKND0 U848 ( .I(port_dest[8]), .ZN(n240) );
  CKND0 U849 ( .I(port_dest[10]), .ZN(n221) );
  AOI33D0 U850 ( .A1(n147), .A2(n358), .A3(n342), .B1(n336), .B2(n87), .B3(
        n355), .ZN(n372) );
  NR2D0 U851 ( .A1(n325), .A2(port_dest[26]), .ZN(n355) );
  CKND0 U852 ( .I(port_dest[25]), .ZN(n87) );
  CKND0 U853 ( .I(port_dest[24]), .ZN(n336) );
  NR2D0 U854 ( .A1(n138), .A2(port_dest[1]), .ZN(n342) );
  CKND0 U855 ( .I(port_dest[3]), .ZN(n138) );
  CKND0 U856 ( .I(port_dest[2]), .ZN(n358) );
  CKND0 U857 ( .I(port_dest[0]), .ZN(n147) );
  AOI33D0 U858 ( .A1(n335), .A2(n107), .A3(n356), .B1(n70), .B2(n48), .B3(n357), .ZN(n371) );
  NR2D0 U859 ( .A1(n50), .A2(port_dest[22]), .ZN(n357) );
  CKND0 U860 ( .I(port_dest[23]), .ZN(n50) );
  CKND0 U861 ( .I(port_dest[21]), .ZN(n48) );
  CKND0 U862 ( .I(port_dest[20]), .ZN(n70) );
  NR2D0 U863 ( .A1(n111), .A2(port_dest[30]), .ZN(n356) );
  CKND0 U864 ( .I(port_dest[29]), .ZN(n107) );
  CKND0 U865 ( .I(port_dest[28]), .ZN(n335) );
  CKND0 U866 ( .I(port_dest[31]), .ZN(n111) );
  CKND0 U867 ( .I(port_dest[27]), .ZN(n325) );
endmodule


module layer_controller ( data_in, data_out, layer_data_in, layer_data_out, 
        addr, len, WE, RE, op_done, rst, layer_en, clk, layer_done );
  input [127:0] data_in;
  output [127:0] data_out;
  input [159:0] layer_data_in;
  output [159:0] layer_data_out;
  output [15:0] addr;
  output [3:0] len;
  input op_done, rst, layer_en, clk;
  output WE, RE, layer_done;
  wire   RE, \input_value[7][127] , \input_value[7][126] ,
         \input_value[7][125] , \input_value[7][124] , \input_value[7][123] ,
         \input_value[7][122] , \input_value[7][121] , \input_value[7][120] ,
         \input_value[7][119] , \input_value[7][118] , \input_value[7][117] ,
         \input_value[7][116] , \input_value[7][115] , \input_value[7][114] ,
         \input_value[7][113] , \input_value[7][112] , \input_value[7][111] ,
         \input_value[7][110] , \input_value[7][109] , \input_value[7][108] ,
         \input_value[7][107] , \input_value[7][106] , \input_value[7][105] ,
         \input_value[7][104] , \input_value[7][103] , \input_value[7][102] ,
         \input_value[7][101] , \input_value[7][100] , \input_value[7][99] ,
         \input_value[7][98] , \input_value[7][97] , \input_value[7][96] ,
         \input_value[7][95] , \input_value[7][94] , \input_value[7][93] ,
         \input_value[7][92] , \input_value[7][91] , \input_value[7][90] ,
         \input_value[7][89] , \input_value[7][88] , \input_value[7][87] ,
         \input_value[7][86] , \input_value[7][85] , \input_value[7][84] ,
         \input_value[7][83] , \input_value[7][82] , \input_value[7][81] ,
         \input_value[7][80] , \input_value[7][79] , \input_value[7][78] ,
         \input_value[7][77] , \input_value[7][76] , \input_value[7][75] ,
         \input_value[7][74] , \input_value[7][73] , \input_value[7][72] ,
         \input_value[7][71] , \input_value[7][70] , \input_value[7][69] ,
         \input_value[7][68] , \input_value[7][67] , \input_value[7][66] ,
         \input_value[7][65] , \input_value[7][64] , \input_value[7][63] ,
         \input_value[7][62] , \input_value[7][61] , \input_value[7][60] ,
         \input_value[7][59] , \input_value[7][58] , \input_value[7][57] ,
         \input_value[7][56] , \input_value[7][55] , \input_value[7][54] ,
         \input_value[7][53] , \input_value[7][52] , \input_value[7][51] ,
         \input_value[7][50] , \input_value[7][49] , \input_value[7][48] ,
         \input_value[7][47] , \input_value[7][46] , \input_value[7][45] ,
         \input_value[7][44] , \input_value[7][43] , \input_value[7][42] ,
         \input_value[7][41] , \input_value[7][40] , \input_value[7][39] ,
         \input_value[7][38] , \input_value[7][37] , \input_value[7][36] ,
         \input_value[7][35] , \input_value[7][34] , \input_value[7][33] ,
         \input_value[7][32] , \input_value[7][31] , \input_value[7][30] ,
         \input_value[7][29] , \input_value[7][28] , \input_value[7][27] ,
         \input_value[7][26] , \input_value[7][25] , \input_value[7][24] ,
         \input_value[7][23] , \input_value[7][22] , \input_value[7][21] ,
         \input_value[7][20] , \input_value[7][19] , \input_value[7][18] ,
         \input_value[7][17] , \input_value[7][16] , \input_value[7][15] ,
         \input_value[7][14] , \input_value[7][13] , \input_value[7][12] ,
         \input_value[7][11] , \input_value[7][10] , \input_value[7][9] ,
         \input_value[7][8] , \input_value[7][7] , \input_value[7][6] ,
         \input_value[7][5] , \input_value[7][4] , \input_value[7][3] ,
         \input_value[7][2] , \input_value[7][1] , \input_value[7][0] ,
         \input_value[6][127] , \input_value[6][126] , \input_value[6][125] ,
         \input_value[6][124] , \input_value[6][123] , \input_value[6][122] ,
         \input_value[6][121] , \input_value[6][120] , \input_value[6][119] ,
         \input_value[6][118] , \input_value[6][117] , \input_value[6][116] ,
         \input_value[6][115] , \input_value[6][114] , \input_value[6][113] ,
         \input_value[6][112] , \input_value[6][111] , \input_value[6][110] ,
         \input_value[6][109] , \input_value[6][108] , \input_value[6][107] ,
         \input_value[6][106] , \input_value[6][105] , \input_value[6][104] ,
         \input_value[6][103] , \input_value[6][102] , \input_value[6][101] ,
         \input_value[6][100] , \input_value[6][99] , \input_value[6][98] ,
         \input_value[6][97] , \input_value[6][96] , \input_value[6][95] ,
         \input_value[6][94] , \input_value[6][93] , \input_value[6][92] ,
         \input_value[6][91] , \input_value[6][90] , \input_value[6][89] ,
         \input_value[6][88] , \input_value[6][87] , \input_value[6][86] ,
         \input_value[6][85] , \input_value[6][84] , \input_value[6][83] ,
         \input_value[6][82] , \input_value[6][81] , \input_value[6][80] ,
         \input_value[6][79] , \input_value[6][78] , \input_value[6][77] ,
         \input_value[6][76] , \input_value[6][75] , \input_value[6][74] ,
         \input_value[6][73] , \input_value[6][72] , \input_value[6][71] ,
         \input_value[6][70] , \input_value[6][69] , \input_value[6][68] ,
         \input_value[6][67] , \input_value[6][66] , \input_value[6][65] ,
         \input_value[6][64] , \input_value[6][63] , \input_value[6][62] ,
         \input_value[6][61] , \input_value[6][60] , \input_value[6][59] ,
         \input_value[6][58] , \input_value[6][57] , \input_value[6][56] ,
         \input_value[6][55] , \input_value[6][54] , \input_value[6][53] ,
         \input_value[6][52] , \input_value[6][51] , \input_value[6][50] ,
         \input_value[6][49] , \input_value[6][48] , \input_value[6][47] ,
         \input_value[6][46] , \input_value[6][45] , \input_value[6][44] ,
         \input_value[6][43] , \input_value[6][42] , \input_value[6][41] ,
         \input_value[6][40] , \input_value[6][39] , \input_value[6][38] ,
         \input_value[6][37] , \input_value[6][36] , \input_value[6][35] ,
         \input_value[6][34] , \input_value[6][33] , \input_value[6][32] ,
         \input_value[6][31] , \input_value[6][30] , \input_value[6][29] ,
         \input_value[6][28] , \input_value[6][27] , \input_value[6][26] ,
         \input_value[6][25] , \input_value[6][24] , \input_value[6][23] ,
         \input_value[6][22] , \input_value[6][21] , \input_value[6][20] ,
         \input_value[6][19] , \input_value[6][18] , \input_value[6][17] ,
         \input_value[6][16] , \input_value[6][15] , \input_value[6][14] ,
         \input_value[6][13] , \input_value[6][12] , \input_value[6][11] ,
         \input_value[6][10] , \input_value[6][9] , \input_value[6][8] ,
         \input_value[6][7] , \input_value[6][6] , \input_value[6][5] ,
         \input_value[6][4] , \input_value[6][3] , \input_value[6][2] ,
         \input_value[6][1] , \input_value[6][0] , \input_value[5][127] ,
         \input_value[5][126] , \input_value[5][125] , \input_value[5][124] ,
         \input_value[5][123] , \input_value[5][122] , \input_value[5][121] ,
         \input_value[5][120] , \input_value[5][119] , \input_value[5][118] ,
         \input_value[5][117] , \input_value[5][116] , \input_value[5][115] ,
         \input_value[5][114] , \input_value[5][113] , \input_value[5][112] ,
         \input_value[5][111] , \input_value[5][110] , \input_value[5][109] ,
         \input_value[5][108] , \input_value[5][107] , \input_value[5][106] ,
         \input_value[5][105] , \input_value[5][104] , \input_value[5][103] ,
         \input_value[5][102] , \input_value[5][101] , \input_value[5][100] ,
         \input_value[5][99] , \input_value[5][98] , \input_value[5][97] ,
         \input_value[5][96] , \input_value[5][95] , \input_value[5][94] ,
         \input_value[5][93] , \input_value[5][92] , \input_value[5][91] ,
         \input_value[5][90] , \input_value[5][89] , \input_value[5][88] ,
         \input_value[5][87] , \input_value[5][86] , \input_value[5][85] ,
         \input_value[5][84] , \input_value[5][83] , \input_value[5][82] ,
         \input_value[5][81] , \input_value[5][80] , \input_value[5][79] ,
         \input_value[5][78] , \input_value[5][77] , \input_value[5][76] ,
         \input_value[5][75] , \input_value[5][74] , \input_value[5][73] ,
         \input_value[5][72] , \input_value[5][71] , \input_value[5][70] ,
         \input_value[5][69] , \input_value[5][68] , \input_value[5][67] ,
         \input_value[5][66] , \input_value[5][65] , \input_value[5][64] ,
         \input_value[5][63] , \input_value[5][62] , \input_value[5][61] ,
         \input_value[5][60] , \input_value[5][59] , \input_value[5][58] ,
         \input_value[5][57] , \input_value[5][56] , \input_value[5][55] ,
         \input_value[5][54] , \input_value[5][53] , \input_value[5][52] ,
         \input_value[5][51] , \input_value[5][50] , \input_value[5][49] ,
         \input_value[5][48] , \input_value[5][47] , \input_value[5][46] ,
         \input_value[5][45] , \input_value[5][44] , \input_value[5][43] ,
         \input_value[5][42] , \input_value[5][41] , \input_value[5][40] ,
         \input_value[5][39] , \input_value[5][38] , \input_value[5][37] ,
         \input_value[5][36] , \input_value[5][35] , \input_value[5][34] ,
         \input_value[5][33] , \input_value[5][32] , \input_value[5][31] ,
         \input_value[5][30] , \input_value[5][29] , \input_value[5][28] ,
         \input_value[5][27] , \input_value[5][26] , \input_value[5][25] ,
         \input_value[5][24] , \input_value[5][23] , \input_value[5][22] ,
         \input_value[5][21] , \input_value[5][20] , \input_value[5][19] ,
         \input_value[5][18] , \input_value[5][17] , \input_value[5][16] ,
         \input_value[5][15] , \input_value[5][14] , \input_value[5][13] ,
         \input_value[5][12] , \input_value[5][11] , \input_value[5][10] ,
         \input_value[5][9] , \input_value[5][8] , \input_value[5][7] ,
         \input_value[5][6] , \input_value[5][5] , \input_value[5][4] ,
         \input_value[5][3] , \input_value[5][2] , \input_value[5][1] ,
         \input_value[5][0] , \input_value[4][127] , \input_value[4][126] ,
         \input_value[4][125] , \input_value[4][124] , \input_value[4][123] ,
         \input_value[4][122] , \input_value[4][121] , \input_value[4][120] ,
         \input_value[4][119] , \input_value[4][118] , \input_value[4][117] ,
         \input_value[4][116] , \input_value[4][115] , \input_value[4][114] ,
         \input_value[4][113] , \input_value[4][112] , \input_value[4][111] ,
         \input_value[4][110] , \input_value[4][109] , \input_value[4][108] ,
         \input_value[4][107] , \input_value[4][106] , \input_value[4][105] ,
         \input_value[4][104] , \input_value[4][103] , \input_value[4][102] ,
         \input_value[4][101] , \input_value[4][100] , \input_value[4][99] ,
         \input_value[4][98] , \input_value[4][97] , \input_value[4][96] ,
         \input_value[4][95] , \input_value[4][94] , \input_value[4][93] ,
         \input_value[4][92] , \input_value[4][91] , \input_value[4][90] ,
         \input_value[4][89] , \input_value[4][88] , \input_value[4][87] ,
         \input_value[4][86] , \input_value[4][85] , \input_value[4][84] ,
         \input_value[4][83] , \input_value[4][82] , \input_value[4][81] ,
         \input_value[4][80] , \input_value[4][79] , \input_value[4][78] ,
         \input_value[4][77] , \input_value[4][76] , \input_value[4][75] ,
         \input_value[4][74] , \input_value[4][73] , \input_value[4][72] ,
         \input_value[4][71] , \input_value[4][70] , \input_value[4][69] ,
         \input_value[4][68] , \input_value[4][67] , \input_value[4][66] ,
         \input_value[4][65] , \input_value[4][64] , \input_value[4][63] ,
         \input_value[4][62] , \input_value[4][61] , \input_value[4][60] ,
         \input_value[4][59] , \input_value[4][58] , \input_value[4][57] ,
         \input_value[4][56] , \input_value[4][55] , \input_value[4][54] ,
         \input_value[4][53] , \input_value[4][52] , \input_value[4][51] ,
         \input_value[4][50] , \input_value[4][49] , \input_value[4][48] ,
         \input_value[4][47] , \input_value[4][46] , \input_value[4][45] ,
         \input_value[4][44] , \input_value[4][43] , \input_value[4][42] ,
         \input_value[4][41] , \input_value[4][40] , \input_value[4][39] ,
         \input_value[4][38] , \input_value[4][37] , \input_value[4][36] ,
         \input_value[4][35] , \input_value[4][34] , \input_value[4][33] ,
         \input_value[4][32] , \input_value[4][31] , \input_value[4][30] ,
         \input_value[4][29] , \input_value[4][28] , \input_value[4][27] ,
         \input_value[4][26] , \input_value[4][25] , \input_value[4][24] ,
         \input_value[4][23] , \input_value[4][22] , \input_value[4][21] ,
         \input_value[4][20] , \input_value[4][19] , \input_value[4][18] ,
         \input_value[4][17] , \input_value[4][16] , \input_value[4][15] ,
         \input_value[4][14] , \input_value[4][13] , \input_value[4][12] ,
         \input_value[4][11] , \input_value[4][10] , \input_value[4][9] ,
         \input_value[4][8] , \input_value[4][7] , \input_value[4][6] ,
         \input_value[4][5] , \input_value[4][4] , \input_value[4][3] ,
         \input_value[4][2] , \input_value[4][1] , \input_value[4][0] ,
         \input_value[3][127] , \input_value[3][126] , \input_value[3][125] ,
         \input_value[3][124] , \input_value[3][123] , \input_value[3][122] ,
         \input_value[3][121] , \input_value[3][120] , \input_value[3][119] ,
         \input_value[3][118] , \input_value[3][117] , \input_value[3][116] ,
         \input_value[3][115] , \input_value[3][114] , \input_value[3][113] ,
         \input_value[3][112] , \input_value[3][111] , \input_value[3][110] ,
         \input_value[3][109] , \input_value[3][108] , \input_value[3][107] ,
         \input_value[3][106] , \input_value[3][105] , \input_value[3][104] ,
         \input_value[3][103] , \input_value[3][102] , \input_value[3][101] ,
         \input_value[3][100] , \input_value[3][99] , \input_value[3][98] ,
         \input_value[3][97] , \input_value[3][96] , \input_value[3][95] ,
         \input_value[3][94] , \input_value[3][93] , \input_value[3][92] ,
         \input_value[3][91] , \input_value[3][90] , \input_value[3][89] ,
         \input_value[3][88] , \input_value[3][87] , \input_value[3][86] ,
         \input_value[3][85] , \input_value[3][84] , \input_value[3][83] ,
         \input_value[3][82] , \input_value[3][81] , \input_value[3][80] ,
         \input_value[3][79] , \input_value[3][78] , \input_value[3][77] ,
         \input_value[3][76] , \input_value[3][75] , \input_value[3][74] ,
         \input_value[3][73] , \input_value[3][72] , \input_value[3][71] ,
         \input_value[3][70] , \input_value[3][69] , \input_value[3][68] ,
         \input_value[3][67] , \input_value[3][66] , \input_value[3][65] ,
         \input_value[3][64] , \input_value[3][63] , \input_value[3][62] ,
         \input_value[3][61] , \input_value[3][60] , \input_value[3][59] ,
         \input_value[3][58] , \input_value[3][57] , \input_value[3][56] ,
         \input_value[3][55] , \input_value[3][54] , \input_value[3][53] ,
         \input_value[3][52] , \input_value[3][51] , \input_value[3][50] ,
         \input_value[3][49] , \input_value[3][48] , \input_value[3][47] ,
         \input_value[3][46] , \input_value[3][45] , \input_value[3][44] ,
         \input_value[3][43] , \input_value[3][42] , \input_value[3][41] ,
         \input_value[3][40] , \input_value[3][39] , \input_value[3][38] ,
         \input_value[3][37] , \input_value[3][36] , \input_value[3][35] ,
         \input_value[3][34] , \input_value[3][33] , \input_value[3][32] ,
         \input_value[3][31] , \input_value[3][30] , \input_value[3][29] ,
         \input_value[3][28] , \input_value[3][27] , \input_value[3][26] ,
         \input_value[3][25] , \input_value[3][24] , \input_value[3][23] ,
         \input_value[3][22] , \input_value[3][21] , \input_value[3][20] ,
         \input_value[3][19] , \input_value[3][18] , \input_value[3][17] ,
         \input_value[3][16] , \input_value[3][15] , \input_value[3][14] ,
         \input_value[3][13] , \input_value[3][12] , \input_value[3][11] ,
         \input_value[3][10] , \input_value[3][9] , \input_value[3][8] ,
         \input_value[3][7] , \input_value[3][6] , \input_value[3][5] ,
         \input_value[3][4] , \input_value[3][3] , \input_value[3][2] ,
         \input_value[3][1] , \input_value[3][0] , \input_value[2][127] ,
         \input_value[2][126] , \input_value[2][125] , \input_value[2][124] ,
         \input_value[2][123] , \input_value[2][122] , \input_value[2][121] ,
         \input_value[2][120] , \input_value[2][119] , \input_value[2][118] ,
         \input_value[2][117] , \input_value[2][116] , \input_value[2][115] ,
         \input_value[2][114] , \input_value[2][113] , \input_value[2][112] ,
         \input_value[2][111] , \input_value[2][110] , \input_value[2][109] ,
         \input_value[2][108] , \input_value[2][107] , \input_value[2][106] ,
         \input_value[2][105] , \input_value[2][104] , \input_value[2][103] ,
         \input_value[2][102] , \input_value[2][101] , \input_value[2][100] ,
         \input_value[2][99] , \input_value[2][98] , \input_value[2][97] ,
         \input_value[2][96] , \input_value[2][95] , \input_value[2][94] ,
         \input_value[2][93] , \input_value[2][92] , \input_value[2][91] ,
         \input_value[2][90] , \input_value[2][89] , \input_value[2][88] ,
         \input_value[2][87] , \input_value[2][86] , \input_value[2][85] ,
         \input_value[2][84] , \input_value[2][83] , \input_value[2][82] ,
         \input_value[2][81] , \input_value[2][80] , \input_value[2][79] ,
         \input_value[2][78] , \input_value[2][77] , \input_value[2][76] ,
         \input_value[2][75] , \input_value[2][74] , \input_value[2][73] ,
         \input_value[2][72] , \input_value[2][71] , \input_value[2][70] ,
         \input_value[2][69] , \input_value[2][68] , \input_value[2][67] ,
         \input_value[2][66] , \input_value[2][65] , \input_value[2][64] ,
         \input_value[2][63] , \input_value[2][62] , \input_value[2][61] ,
         \input_value[2][60] , \input_value[2][59] , \input_value[2][58] ,
         \input_value[2][57] , \input_value[2][56] , \input_value[2][55] ,
         \input_value[2][54] , \input_value[2][53] , \input_value[2][52] ,
         \input_value[2][51] , \input_value[2][50] , \input_value[2][49] ,
         \input_value[2][48] , \input_value[2][47] , \input_value[2][46] ,
         \input_value[2][45] , \input_value[2][44] , \input_value[2][43] ,
         \input_value[2][42] , \input_value[2][41] , \input_value[2][40] ,
         \input_value[2][39] , \input_value[2][38] , \input_value[2][37] ,
         \input_value[2][36] , \input_value[2][35] , \input_value[2][34] ,
         \input_value[2][33] , \input_value[2][32] , \input_value[2][31] ,
         \input_value[2][30] , \input_value[2][29] , \input_value[2][28] ,
         \input_value[2][27] , \input_value[2][26] , \input_value[2][25] ,
         \input_value[2][24] , \input_value[2][23] , \input_value[2][22] ,
         \input_value[2][21] , \input_value[2][20] , \input_value[2][19] ,
         \input_value[2][18] , \input_value[2][17] , \input_value[2][16] ,
         \input_value[2][15] , \input_value[2][14] , \input_value[2][13] ,
         \input_value[2][12] , \input_value[2][11] , \input_value[2][10] ,
         \input_value[2][9] , \input_value[2][8] , \input_value[2][7] ,
         \input_value[2][6] , \input_value[2][5] , \input_value[2][4] ,
         \input_value[2][3] , \input_value[2][2] , \input_value[2][1] ,
         \input_value[2][0] , \input_value[1][127] , \input_value[1][126] ,
         \input_value[1][125] , \input_value[1][124] , \input_value[1][123] ,
         \input_value[1][122] , \input_value[1][121] , \input_value[1][120] ,
         \input_value[1][119] , \input_value[1][118] , \input_value[1][117] ,
         \input_value[1][116] , \input_value[1][115] , \input_value[1][114] ,
         \input_value[1][113] , \input_value[1][112] , \input_value[1][111] ,
         \input_value[1][110] , \input_value[1][109] , \input_value[1][108] ,
         \input_value[1][107] , \input_value[1][106] , \input_value[1][105] ,
         \input_value[1][104] , \input_value[1][103] , \input_value[1][102] ,
         \input_value[1][101] , \input_value[1][100] , \input_value[1][99] ,
         \input_value[1][98] , \input_value[1][97] , \input_value[1][96] ,
         \input_value[1][95] , \input_value[1][94] , \input_value[1][93] ,
         \input_value[1][92] , \input_value[1][91] , \input_value[1][90] ,
         \input_value[1][89] , \input_value[1][88] , \input_value[1][87] ,
         \input_value[1][86] , \input_value[1][85] , \input_value[1][84] ,
         \input_value[1][83] , \input_value[1][82] , \input_value[1][81] ,
         \input_value[1][80] , \input_value[1][79] , \input_value[1][78] ,
         \input_value[1][77] , \input_value[1][76] , \input_value[1][75] ,
         \input_value[1][74] , \input_value[1][73] , \input_value[1][72] ,
         \input_value[1][71] , \input_value[1][70] , \input_value[1][69] ,
         \input_value[1][68] , \input_value[1][67] , \input_value[1][66] ,
         \input_value[1][65] , \input_value[1][64] , \input_value[1][63] ,
         \input_value[1][62] , \input_value[1][61] , \input_value[1][60] ,
         \input_value[1][59] , \input_value[1][58] , \input_value[1][57] ,
         \input_value[1][56] , \input_value[1][55] , \input_value[1][54] ,
         \input_value[1][53] , \input_value[1][52] , \input_value[1][51] ,
         \input_value[1][50] , \input_value[1][49] , \input_value[1][48] ,
         \input_value[1][47] , \input_value[1][46] , \input_value[1][45] ,
         \input_value[1][44] , \input_value[1][43] , \input_value[1][42] ,
         \input_value[1][41] , \input_value[1][40] , \input_value[1][39] ,
         \input_value[1][38] , \input_value[1][37] , \input_value[1][36] ,
         \input_value[1][35] , \input_value[1][34] , \input_value[1][33] ,
         \input_value[1][32] , \input_value[1][31] , \input_value[1][30] ,
         \input_value[1][29] , \input_value[1][28] , \input_value[1][27] ,
         \input_value[1][26] , \input_value[1][25] , \input_value[1][24] ,
         \input_value[1][23] , \input_value[1][22] , \input_value[1][21] ,
         \input_value[1][20] , \input_value[1][19] , \input_value[1][18] ,
         \input_value[1][17] , \input_value[1][16] , \input_value[1][15] ,
         \input_value[1][14] , \input_value[1][13] , \input_value[1][12] ,
         \input_value[1][11] , \input_value[1][10] , \input_value[1][9] ,
         \input_value[1][8] , \input_value[1][7] , \input_value[1][6] ,
         \input_value[1][5] , \input_value[1][4] , \input_value[1][3] ,
         \input_value[1][2] , \input_value[1][1] , \input_value[1][0] ,
         \input_value[0][127] , \input_value[0][126] , \input_value[0][125] ,
         \input_value[0][124] , \input_value[0][123] , \input_value[0][122] ,
         \input_value[0][121] , \input_value[0][120] , \input_value[0][119] ,
         \input_value[0][118] , \input_value[0][117] , \input_value[0][116] ,
         \input_value[0][115] , \input_value[0][114] , \input_value[0][113] ,
         \input_value[0][112] , \input_value[0][111] , \input_value[0][110] ,
         \input_value[0][109] , \input_value[0][108] , \input_value[0][107] ,
         \input_value[0][106] , \input_value[0][105] , \input_value[0][104] ,
         \input_value[0][103] , \input_value[0][102] , \input_value[0][101] ,
         \input_value[0][100] , \input_value[0][99] , \input_value[0][98] ,
         \input_value[0][97] , \input_value[0][96] , \input_value[0][95] ,
         \input_value[0][94] , \input_value[0][93] , \input_value[0][92] ,
         \input_value[0][91] , \input_value[0][90] , \input_value[0][89] ,
         \input_value[0][88] , \input_value[0][87] , \input_value[0][86] ,
         \input_value[0][85] , \input_value[0][84] , \input_value[0][83] ,
         \input_value[0][82] , \input_value[0][81] , \input_value[0][80] ,
         \input_value[0][79] , \input_value[0][78] , \input_value[0][77] ,
         \input_value[0][76] , \input_value[0][75] , \input_value[0][74] ,
         \input_value[0][73] , \input_value[0][72] , \input_value[0][71] ,
         \input_value[0][70] , \input_value[0][69] , \input_value[0][68] ,
         \input_value[0][67] , \input_value[0][66] , \input_value[0][65] ,
         \input_value[0][64] , \input_value[0][63] , \input_value[0][62] ,
         \input_value[0][61] , \input_value[0][60] , \input_value[0][59] ,
         \input_value[0][58] , \input_value[0][57] , \input_value[0][56] ,
         \input_value[0][55] , \input_value[0][54] , \input_value[0][53] ,
         \input_value[0][52] , \input_value[0][51] , \input_value[0][50] ,
         \input_value[0][49] , \input_value[0][48] , \input_value[0][47] ,
         \input_value[0][46] , \input_value[0][45] , \input_value[0][44] ,
         \input_value[0][43] , \input_value[0][42] , \input_value[0][41] ,
         \input_value[0][40] , \input_value[0][39] , \input_value[0][38] ,
         \input_value[0][37] , \input_value[0][36] , \input_value[0][35] ,
         \input_value[0][34] , \input_value[0][33] , \input_value[0][32] ,
         \input_value[0][31] , \input_value[0][30] , \input_value[0][29] ,
         \input_value[0][28] , \input_value[0][27] , \input_value[0][26] ,
         \input_value[0][25] , \input_value[0][24] , \input_value[0][23] ,
         \input_value[0][22] , \input_value[0][21] , \input_value[0][20] ,
         \input_value[0][19] , \input_value[0][18] , \input_value[0][17] ,
         \input_value[0][16] , \input_value[0][15] , \input_value[0][14] ,
         \input_value[0][13] , \input_value[0][12] , \input_value[0][11] ,
         \input_value[0][10] , \input_value[0][9] , \input_value[0][8] ,
         \input_value[0][7] , \input_value[0][6] , \input_value[0][5] ,
         \input_value[0][4] , \input_value[0][3] , \input_value[0][2] ,
         \input_value[0][1] , \input_value[0][0] , \input_weight[7][127] ,
         \input_weight[7][126] , \input_weight[7][125] ,
         \input_weight[7][124] , \input_weight[7][123] ,
         \input_weight[7][122] , \input_weight[7][121] ,
         \input_weight[7][120] , \input_weight[7][119] ,
         \input_weight[7][118] , \input_weight[7][117] ,
         \input_weight[7][116] , \input_weight[7][115] ,
         \input_weight[7][114] , \input_weight[7][113] ,
         \input_weight[7][112] , \input_weight[7][111] ,
         \input_weight[7][110] , \input_weight[7][109] ,
         \input_weight[7][108] , \input_weight[7][107] ,
         \input_weight[7][106] , \input_weight[7][105] ,
         \input_weight[7][104] , \input_weight[7][103] ,
         \input_weight[7][102] , \input_weight[7][101] ,
         \input_weight[7][100] , \input_weight[7][99] , \input_weight[7][98] ,
         \input_weight[7][97] , \input_weight[7][96] , \input_weight[7][95] ,
         \input_weight[7][94] , \input_weight[7][93] , \input_weight[7][92] ,
         \input_weight[7][91] , \input_weight[7][90] , \input_weight[7][89] ,
         \input_weight[7][88] , \input_weight[7][87] , \input_weight[7][86] ,
         \input_weight[7][85] , \input_weight[7][84] , \input_weight[7][83] ,
         \input_weight[7][82] , \input_weight[7][81] , \input_weight[7][80] ,
         \input_weight[7][79] , \input_weight[7][78] , \input_weight[7][77] ,
         \input_weight[7][76] , \input_weight[7][75] , \input_weight[7][74] ,
         \input_weight[7][73] , \input_weight[7][72] , \input_weight[7][71] ,
         \input_weight[7][70] , \input_weight[7][69] , \input_weight[7][68] ,
         \input_weight[7][67] , \input_weight[7][66] , \input_weight[7][65] ,
         \input_weight[7][64] , \input_weight[7][63] , \input_weight[7][62] ,
         \input_weight[7][61] , \input_weight[7][60] , \input_weight[7][59] ,
         \input_weight[7][58] , \input_weight[7][57] , \input_weight[7][56] ,
         \input_weight[7][55] , \input_weight[7][54] , \input_weight[7][53] ,
         \input_weight[7][52] , \input_weight[7][51] , \input_weight[7][50] ,
         \input_weight[7][49] , \input_weight[7][48] , \input_weight[7][47] ,
         \input_weight[7][46] , \input_weight[7][45] , \input_weight[7][44] ,
         \input_weight[7][43] , \input_weight[7][42] , \input_weight[7][41] ,
         \input_weight[7][40] , \input_weight[7][39] , \input_weight[7][38] ,
         \input_weight[7][37] , \input_weight[7][36] , \input_weight[7][35] ,
         \input_weight[7][34] , \input_weight[7][33] , \input_weight[7][32] ,
         \input_weight[7][31] , \input_weight[7][30] , \input_weight[7][29] ,
         \input_weight[7][28] , \input_weight[7][27] , \input_weight[7][26] ,
         \input_weight[7][25] , \input_weight[7][24] , \input_weight[7][23] ,
         \input_weight[7][22] , \input_weight[7][21] , \input_weight[7][20] ,
         \input_weight[7][19] , \input_weight[7][18] , \input_weight[7][17] ,
         \input_weight[7][16] , \input_weight[7][15] , \input_weight[7][14] ,
         \input_weight[7][13] , \input_weight[7][12] , \input_weight[7][11] ,
         \input_weight[7][10] , \input_weight[7][9] , \input_weight[7][8] ,
         \input_weight[7][7] , \input_weight[7][6] , \input_weight[7][5] ,
         \input_weight[7][4] , \input_weight[7][3] , \input_weight[7][2] ,
         \input_weight[7][1] , \input_weight[7][0] , \input_weight[6][127] ,
         \input_weight[6][126] , \input_weight[6][125] ,
         \input_weight[6][124] , \input_weight[6][123] ,
         \input_weight[6][122] , \input_weight[6][121] ,
         \input_weight[6][120] , \input_weight[6][119] ,
         \input_weight[6][118] , \input_weight[6][117] ,
         \input_weight[6][116] , \input_weight[6][115] ,
         \input_weight[6][114] , \input_weight[6][113] ,
         \input_weight[6][112] , \input_weight[6][111] ,
         \input_weight[6][110] , \input_weight[6][109] ,
         \input_weight[6][108] , \input_weight[6][107] ,
         \input_weight[6][106] , \input_weight[6][105] ,
         \input_weight[6][104] , \input_weight[6][103] ,
         \input_weight[6][102] , \input_weight[6][101] ,
         \input_weight[6][100] , \input_weight[6][99] , \input_weight[6][98] ,
         \input_weight[6][97] , \input_weight[6][96] , \input_weight[6][95] ,
         \input_weight[6][94] , \input_weight[6][93] , \input_weight[6][92] ,
         \input_weight[6][91] , \input_weight[6][90] , \input_weight[6][89] ,
         \input_weight[6][88] , \input_weight[6][87] , \input_weight[6][86] ,
         \input_weight[6][85] , \input_weight[6][84] , \input_weight[6][83] ,
         \input_weight[6][82] , \input_weight[6][81] , \input_weight[6][80] ,
         \input_weight[6][79] , \input_weight[6][78] , \input_weight[6][77] ,
         \input_weight[6][76] , \input_weight[6][75] , \input_weight[6][74] ,
         \input_weight[6][73] , \input_weight[6][72] , \input_weight[6][71] ,
         \input_weight[6][70] , \input_weight[6][69] , \input_weight[6][68] ,
         \input_weight[6][67] , \input_weight[6][66] , \input_weight[6][65] ,
         \input_weight[6][64] , \input_weight[6][63] , \input_weight[6][62] ,
         \input_weight[6][61] , \input_weight[6][60] , \input_weight[6][59] ,
         \input_weight[6][58] , \input_weight[6][57] , \input_weight[6][56] ,
         \input_weight[6][55] , \input_weight[6][54] , \input_weight[6][53] ,
         \input_weight[6][52] , \input_weight[6][51] , \input_weight[6][50] ,
         \input_weight[6][49] , \input_weight[6][48] , \input_weight[6][47] ,
         \input_weight[6][46] , \input_weight[6][45] , \input_weight[6][44] ,
         \input_weight[6][43] , \input_weight[6][42] , \input_weight[6][41] ,
         \input_weight[6][40] , \input_weight[6][39] , \input_weight[6][38] ,
         \input_weight[6][37] , \input_weight[6][36] , \input_weight[6][35] ,
         \input_weight[6][34] , \input_weight[6][33] , \input_weight[6][32] ,
         \input_weight[6][31] , \input_weight[6][30] , \input_weight[6][29] ,
         \input_weight[6][28] , \input_weight[6][27] , \input_weight[6][26] ,
         \input_weight[6][25] , \input_weight[6][24] , \input_weight[6][23] ,
         \input_weight[6][22] , \input_weight[6][21] , \input_weight[6][20] ,
         \input_weight[6][19] , \input_weight[6][18] , \input_weight[6][17] ,
         \input_weight[6][16] , \input_weight[6][15] , \input_weight[6][14] ,
         \input_weight[6][13] , \input_weight[6][12] , \input_weight[6][11] ,
         \input_weight[6][10] , \input_weight[6][9] , \input_weight[6][8] ,
         \input_weight[6][7] , \input_weight[6][6] , \input_weight[6][5] ,
         \input_weight[6][4] , \input_weight[6][3] , \input_weight[6][2] ,
         \input_weight[6][1] , \input_weight[6][0] , \input_weight[5][127] ,
         \input_weight[5][126] , \input_weight[5][125] ,
         \input_weight[5][124] , \input_weight[5][123] ,
         \input_weight[5][122] , \input_weight[5][121] ,
         \input_weight[5][120] , \input_weight[5][119] ,
         \input_weight[5][118] , \input_weight[5][117] ,
         \input_weight[5][116] , \input_weight[5][115] ,
         \input_weight[5][114] , \input_weight[5][113] ,
         \input_weight[5][112] , \input_weight[5][111] ,
         \input_weight[5][110] , \input_weight[5][109] ,
         \input_weight[5][108] , \input_weight[5][107] ,
         \input_weight[5][106] , \input_weight[5][105] ,
         \input_weight[5][104] , \input_weight[5][103] ,
         \input_weight[5][102] , \input_weight[5][101] ,
         \input_weight[5][100] , \input_weight[5][99] , \input_weight[5][98] ,
         \input_weight[5][97] , \input_weight[5][96] , \input_weight[5][95] ,
         \input_weight[5][94] , \input_weight[5][93] , \input_weight[5][92] ,
         \input_weight[5][91] , \input_weight[5][90] , \input_weight[5][89] ,
         \input_weight[5][88] , \input_weight[5][87] , \input_weight[5][86] ,
         \input_weight[5][85] , \input_weight[5][84] , \input_weight[5][83] ,
         \input_weight[5][82] , \input_weight[5][81] , \input_weight[5][80] ,
         \input_weight[5][79] , \input_weight[5][78] , \input_weight[5][77] ,
         \input_weight[5][76] , \input_weight[5][75] , \input_weight[5][74] ,
         \input_weight[5][73] , \input_weight[5][72] , \input_weight[5][71] ,
         \input_weight[5][70] , \input_weight[5][69] , \input_weight[5][68] ,
         \input_weight[5][67] , \input_weight[5][66] , \input_weight[5][65] ,
         \input_weight[5][64] , \input_weight[5][63] , \input_weight[5][62] ,
         \input_weight[5][61] , \input_weight[5][60] , \input_weight[5][59] ,
         \input_weight[5][58] , \input_weight[5][57] , \input_weight[5][56] ,
         \input_weight[5][55] , \input_weight[5][54] , \input_weight[5][53] ,
         \input_weight[5][52] , \input_weight[5][51] , \input_weight[5][50] ,
         \input_weight[5][49] , \input_weight[5][48] , \input_weight[5][47] ,
         \input_weight[5][46] , \input_weight[5][45] , \input_weight[5][44] ,
         \input_weight[5][43] , \input_weight[5][42] , \input_weight[5][41] ,
         \input_weight[5][40] , \input_weight[5][39] , \input_weight[5][38] ,
         \input_weight[5][37] , \input_weight[5][36] , \input_weight[5][35] ,
         \input_weight[5][34] , \input_weight[5][33] , \input_weight[5][32] ,
         \input_weight[5][31] , \input_weight[5][30] , \input_weight[5][29] ,
         \input_weight[5][28] , \input_weight[5][27] , \input_weight[5][26] ,
         \input_weight[5][25] , \input_weight[5][24] , \input_weight[5][23] ,
         \input_weight[5][22] , \input_weight[5][21] , \input_weight[5][20] ,
         \input_weight[5][19] , \input_weight[5][18] , \input_weight[5][17] ,
         \input_weight[5][16] , \input_weight[5][15] , \input_weight[5][14] ,
         \input_weight[5][13] , \input_weight[5][12] , \input_weight[5][11] ,
         \input_weight[5][10] , \input_weight[5][9] , \input_weight[5][8] ,
         \input_weight[5][7] , \input_weight[5][6] , \input_weight[5][5] ,
         \input_weight[5][4] , \input_weight[5][3] , \input_weight[5][2] ,
         \input_weight[5][1] , \input_weight[5][0] , \input_weight[4][127] ,
         \input_weight[4][126] , \input_weight[4][125] ,
         \input_weight[4][124] , \input_weight[4][123] ,
         \input_weight[4][122] , \input_weight[4][121] ,
         \input_weight[4][120] , \input_weight[4][119] ,
         \input_weight[4][118] , \input_weight[4][117] ,
         \input_weight[4][116] , \input_weight[4][115] ,
         \input_weight[4][114] , \input_weight[4][113] ,
         \input_weight[4][112] , \input_weight[4][111] ,
         \input_weight[4][110] , \input_weight[4][109] ,
         \input_weight[4][108] , \input_weight[4][107] ,
         \input_weight[4][106] , \input_weight[4][105] ,
         \input_weight[4][104] , \input_weight[4][103] ,
         \input_weight[4][102] , \input_weight[4][101] ,
         \input_weight[4][100] , \input_weight[4][99] , \input_weight[4][98] ,
         \input_weight[4][97] , \input_weight[4][96] , \input_weight[4][95] ,
         \input_weight[4][94] , \input_weight[4][93] , \input_weight[4][92] ,
         \input_weight[4][91] , \input_weight[4][90] , \input_weight[4][89] ,
         \input_weight[4][88] , \input_weight[4][87] , \input_weight[4][86] ,
         \input_weight[4][85] , \input_weight[4][84] , \input_weight[4][83] ,
         \input_weight[4][82] , \input_weight[4][81] , \input_weight[4][80] ,
         \input_weight[4][79] , \input_weight[4][78] , \input_weight[4][77] ,
         \input_weight[4][76] , \input_weight[4][75] , \input_weight[4][74] ,
         \input_weight[4][73] , \input_weight[4][72] , \input_weight[4][71] ,
         \input_weight[4][70] , \input_weight[4][69] , \input_weight[4][68] ,
         \input_weight[4][67] , \input_weight[4][66] , \input_weight[4][65] ,
         \input_weight[4][64] , \input_weight[4][63] , \input_weight[4][62] ,
         \input_weight[4][61] , \input_weight[4][60] , \input_weight[4][59] ,
         \input_weight[4][58] , \input_weight[4][57] , \input_weight[4][56] ,
         \input_weight[4][55] , \input_weight[4][54] , \input_weight[4][53] ,
         \input_weight[4][52] , \input_weight[4][51] , \input_weight[4][50] ,
         \input_weight[4][49] , \input_weight[4][48] , \input_weight[4][47] ,
         \input_weight[4][46] , \input_weight[4][45] , \input_weight[4][44] ,
         \input_weight[4][43] , \input_weight[4][42] , \input_weight[4][41] ,
         \input_weight[4][40] , \input_weight[4][39] , \input_weight[4][38] ,
         \input_weight[4][37] , \input_weight[4][36] , \input_weight[4][35] ,
         \input_weight[4][34] , \input_weight[4][33] , \input_weight[4][32] ,
         \input_weight[4][31] , \input_weight[4][30] , \input_weight[4][29] ,
         \input_weight[4][28] , \input_weight[4][27] , \input_weight[4][26] ,
         \input_weight[4][25] , \input_weight[4][24] , \input_weight[4][23] ,
         \input_weight[4][22] , \input_weight[4][21] , \input_weight[4][20] ,
         \input_weight[4][19] , \input_weight[4][18] , \input_weight[4][17] ,
         \input_weight[4][16] , \input_weight[4][15] , \input_weight[4][14] ,
         \input_weight[4][13] , \input_weight[4][12] , \input_weight[4][11] ,
         \input_weight[4][10] , \input_weight[4][9] , \input_weight[4][8] ,
         \input_weight[4][7] , \input_weight[4][6] , \input_weight[4][5] ,
         \input_weight[4][4] , \input_weight[4][3] , \input_weight[4][2] ,
         \input_weight[4][1] , \input_weight[4][0] , \input_weight[3][127] ,
         \input_weight[3][126] , \input_weight[3][125] ,
         \input_weight[3][124] , \input_weight[3][123] ,
         \input_weight[3][122] , \input_weight[3][121] ,
         \input_weight[3][120] , \input_weight[3][119] ,
         \input_weight[3][118] , \input_weight[3][117] ,
         \input_weight[3][116] , \input_weight[3][115] ,
         \input_weight[3][114] , \input_weight[3][113] ,
         \input_weight[3][112] , \input_weight[3][111] ,
         \input_weight[3][110] , \input_weight[3][109] ,
         \input_weight[3][108] , \input_weight[3][107] ,
         \input_weight[3][106] , \input_weight[3][105] ,
         \input_weight[3][104] , \input_weight[3][103] ,
         \input_weight[3][102] , \input_weight[3][101] ,
         \input_weight[3][100] , \input_weight[3][99] , \input_weight[3][98] ,
         \input_weight[3][97] , \input_weight[3][96] , \input_weight[3][95] ,
         \input_weight[3][94] , \input_weight[3][93] , \input_weight[3][92] ,
         \input_weight[3][91] , \input_weight[3][90] , \input_weight[3][89] ,
         \input_weight[3][88] , \input_weight[3][87] , \input_weight[3][86] ,
         \input_weight[3][85] , \input_weight[3][84] , \input_weight[3][83] ,
         \input_weight[3][82] , \input_weight[3][81] , \input_weight[3][80] ,
         \input_weight[3][79] , \input_weight[3][78] , \input_weight[3][77] ,
         \input_weight[3][76] , \input_weight[3][75] , \input_weight[3][74] ,
         \input_weight[3][73] , \input_weight[3][72] , \input_weight[3][71] ,
         \input_weight[3][70] , \input_weight[3][69] , \input_weight[3][68] ,
         \input_weight[3][67] , \input_weight[3][66] , \input_weight[3][65] ,
         \input_weight[3][64] , \input_weight[3][63] , \input_weight[3][62] ,
         \input_weight[3][61] , \input_weight[3][60] , \input_weight[3][59] ,
         \input_weight[3][58] , \input_weight[3][57] , \input_weight[3][56] ,
         \input_weight[3][55] , \input_weight[3][54] , \input_weight[3][53] ,
         \input_weight[3][52] , \input_weight[3][51] , \input_weight[3][50] ,
         \input_weight[3][49] , \input_weight[3][48] , \input_weight[3][47] ,
         \input_weight[3][46] , \input_weight[3][45] , \input_weight[3][44] ,
         \input_weight[3][43] , \input_weight[3][42] , \input_weight[3][41] ,
         \input_weight[3][40] , \input_weight[3][39] , \input_weight[3][38] ,
         \input_weight[3][37] , \input_weight[3][36] , \input_weight[3][35] ,
         \input_weight[3][34] , \input_weight[3][33] , \input_weight[3][32] ,
         \input_weight[3][31] , \input_weight[3][30] , \input_weight[3][29] ,
         \input_weight[3][28] , \input_weight[3][27] , \input_weight[3][26] ,
         \input_weight[3][25] , \input_weight[3][24] , \input_weight[3][23] ,
         \input_weight[3][22] , \input_weight[3][21] , \input_weight[3][20] ,
         \input_weight[3][19] , \input_weight[3][18] , \input_weight[3][17] ,
         \input_weight[3][16] , \input_weight[3][15] , \input_weight[3][14] ,
         \input_weight[3][13] , \input_weight[3][12] , \input_weight[3][11] ,
         \input_weight[3][10] , \input_weight[3][9] , \input_weight[3][8] ,
         \input_weight[3][7] , \input_weight[3][6] , \input_weight[3][5] ,
         \input_weight[3][4] , \input_weight[3][3] , \input_weight[3][2] ,
         \input_weight[3][1] , \input_weight[3][0] , \input_weight[2][127] ,
         \input_weight[2][126] , \input_weight[2][125] ,
         \input_weight[2][124] , \input_weight[2][123] ,
         \input_weight[2][122] , \input_weight[2][121] ,
         \input_weight[2][120] , \input_weight[2][119] ,
         \input_weight[2][118] , \input_weight[2][117] ,
         \input_weight[2][116] , \input_weight[2][115] ,
         \input_weight[2][114] , \input_weight[2][113] ,
         \input_weight[2][112] , \input_weight[2][111] ,
         \input_weight[2][110] , \input_weight[2][109] ,
         \input_weight[2][108] , \input_weight[2][107] ,
         \input_weight[2][106] , \input_weight[2][105] ,
         \input_weight[2][104] , \input_weight[2][103] ,
         \input_weight[2][102] , \input_weight[2][101] ,
         \input_weight[2][100] , \input_weight[2][99] , \input_weight[2][98] ,
         \input_weight[2][97] , \input_weight[2][96] , \input_weight[2][95] ,
         \input_weight[2][94] , \input_weight[2][93] , \input_weight[2][92] ,
         \input_weight[2][91] , \input_weight[2][90] , \input_weight[2][89] ,
         \input_weight[2][88] , \input_weight[2][87] , \input_weight[2][86] ,
         \input_weight[2][85] , \input_weight[2][84] , \input_weight[2][83] ,
         \input_weight[2][82] , \input_weight[2][81] , \input_weight[2][80] ,
         \input_weight[2][79] , \input_weight[2][78] , \input_weight[2][77] ,
         \input_weight[2][76] , \input_weight[2][75] , \input_weight[2][74] ,
         \input_weight[2][73] , \input_weight[2][72] , \input_weight[2][71] ,
         \input_weight[2][70] , \input_weight[2][69] , \input_weight[2][68] ,
         \input_weight[2][67] , \input_weight[2][66] , \input_weight[2][65] ,
         \input_weight[2][64] , \input_weight[2][63] , \input_weight[2][62] ,
         \input_weight[2][61] , \input_weight[2][60] , \input_weight[2][59] ,
         \input_weight[2][58] , \input_weight[2][57] , \input_weight[2][56] ,
         \input_weight[2][55] , \input_weight[2][54] , \input_weight[2][53] ,
         \input_weight[2][52] , \input_weight[2][51] , \input_weight[2][50] ,
         \input_weight[2][49] , \input_weight[2][48] , \input_weight[2][47] ,
         \input_weight[2][46] , \input_weight[2][45] , \input_weight[2][44] ,
         \input_weight[2][43] , \input_weight[2][42] , \input_weight[2][41] ,
         \input_weight[2][40] , \input_weight[2][39] , \input_weight[2][38] ,
         \input_weight[2][37] , \input_weight[2][36] , \input_weight[2][35] ,
         \input_weight[2][34] , \input_weight[2][33] , \input_weight[2][32] ,
         \input_weight[2][31] , \input_weight[2][30] , \input_weight[2][29] ,
         \input_weight[2][28] , \input_weight[2][27] , \input_weight[2][26] ,
         \input_weight[2][25] , \input_weight[2][24] , \input_weight[2][23] ,
         \input_weight[2][22] , \input_weight[2][21] , \input_weight[2][20] ,
         \input_weight[2][19] , \input_weight[2][18] , \input_weight[2][17] ,
         \input_weight[2][16] , \input_weight[2][15] , \input_weight[2][14] ,
         \input_weight[2][13] , \input_weight[2][12] , \input_weight[2][11] ,
         \input_weight[2][10] , \input_weight[2][9] , \input_weight[2][8] ,
         \input_weight[2][7] , \input_weight[2][6] , \input_weight[2][5] ,
         \input_weight[2][4] , \input_weight[2][3] , \input_weight[2][2] ,
         \input_weight[2][1] , \input_weight[2][0] , \input_weight[1][127] ,
         \input_weight[1][126] , \input_weight[1][125] ,
         \input_weight[1][124] , \input_weight[1][123] ,
         \input_weight[1][122] , \input_weight[1][121] ,
         \input_weight[1][120] , \input_weight[1][119] ,
         \input_weight[1][118] , \input_weight[1][117] ,
         \input_weight[1][116] , \input_weight[1][115] ,
         \input_weight[1][114] , \input_weight[1][113] ,
         \input_weight[1][112] , \input_weight[1][111] ,
         \input_weight[1][110] , \input_weight[1][109] ,
         \input_weight[1][108] , \input_weight[1][107] ,
         \input_weight[1][106] , \input_weight[1][105] ,
         \input_weight[1][104] , \input_weight[1][103] ,
         \input_weight[1][102] , \input_weight[1][101] ,
         \input_weight[1][100] , \input_weight[1][99] , \input_weight[1][98] ,
         \input_weight[1][97] , \input_weight[1][96] , \input_weight[1][95] ,
         \input_weight[1][94] , \input_weight[1][93] , \input_weight[1][92] ,
         \input_weight[1][91] , \input_weight[1][90] , \input_weight[1][89] ,
         \input_weight[1][88] , \input_weight[1][87] , \input_weight[1][86] ,
         \input_weight[1][85] , \input_weight[1][84] , \input_weight[1][83] ,
         \input_weight[1][82] , \input_weight[1][81] , \input_weight[1][80] ,
         \input_weight[1][79] , \input_weight[1][78] , \input_weight[1][77] ,
         \input_weight[1][76] , \input_weight[1][75] , \input_weight[1][74] ,
         \input_weight[1][73] , \input_weight[1][72] , \input_weight[1][71] ,
         \input_weight[1][70] , \input_weight[1][69] , \input_weight[1][68] ,
         \input_weight[1][67] , \input_weight[1][66] , \input_weight[1][65] ,
         \input_weight[1][64] , \input_weight[1][63] , \input_weight[1][62] ,
         \input_weight[1][61] , \input_weight[1][60] , \input_weight[1][59] ,
         \input_weight[1][58] , \input_weight[1][57] , \input_weight[1][56] ,
         \input_weight[1][55] , \input_weight[1][54] , \input_weight[1][53] ,
         \input_weight[1][52] , \input_weight[1][51] , \input_weight[1][50] ,
         \input_weight[1][49] , \input_weight[1][48] , \input_weight[1][47] ,
         \input_weight[1][46] , \input_weight[1][45] , \input_weight[1][44] ,
         \input_weight[1][43] , \input_weight[1][42] , \input_weight[1][41] ,
         \input_weight[1][40] , \input_weight[1][39] , \input_weight[1][38] ,
         \input_weight[1][37] , \input_weight[1][36] , \input_weight[1][35] ,
         \input_weight[1][34] , \input_weight[1][33] , \input_weight[1][32] ,
         \input_weight[1][31] , \input_weight[1][30] , \input_weight[1][29] ,
         \input_weight[1][28] , \input_weight[1][27] , \input_weight[1][26] ,
         \input_weight[1][25] , \input_weight[1][24] , \input_weight[1][23] ,
         \input_weight[1][22] , \input_weight[1][21] , \input_weight[1][20] ,
         \input_weight[1][19] , \input_weight[1][18] , \input_weight[1][17] ,
         \input_weight[1][16] , \input_weight[1][15] , \input_weight[1][14] ,
         \input_weight[1][13] , \input_weight[1][12] , \input_weight[1][11] ,
         \input_weight[1][10] , \input_weight[1][9] , \input_weight[1][8] ,
         \input_weight[1][7] , \input_weight[1][6] , \input_weight[1][5] ,
         \input_weight[1][4] , \input_weight[1][3] , \input_weight[1][2] ,
         \input_weight[1][1] , \input_weight[1][0] , \input_weight[0][127] ,
         \input_weight[0][126] , \input_weight[0][125] ,
         \input_weight[0][124] , \input_weight[0][123] ,
         \input_weight[0][122] , \input_weight[0][121] ,
         \input_weight[0][120] , \input_weight[0][119] ,
         \input_weight[0][118] , \input_weight[0][117] ,
         \input_weight[0][116] , \input_weight[0][115] ,
         \input_weight[0][114] , \input_weight[0][113] ,
         \input_weight[0][112] , \input_weight[0][111] ,
         \input_weight[0][110] , \input_weight[0][109] ,
         \input_weight[0][108] , \input_weight[0][107] ,
         \input_weight[0][106] , \input_weight[0][105] ,
         \input_weight[0][104] , \input_weight[0][103] ,
         \input_weight[0][102] , \input_weight[0][101] ,
         \input_weight[0][100] , \input_weight[0][99] , \input_weight[0][98] ,
         \input_weight[0][97] , \input_weight[0][96] , \input_weight[0][95] ,
         \input_weight[0][94] , \input_weight[0][93] , \input_weight[0][92] ,
         \input_weight[0][91] , \input_weight[0][90] , \input_weight[0][89] ,
         \input_weight[0][88] , \input_weight[0][87] , \input_weight[0][86] ,
         \input_weight[0][85] , \input_weight[0][84] , \input_weight[0][83] ,
         \input_weight[0][82] , \input_weight[0][81] , \input_weight[0][80] ,
         \input_weight[0][79] , \input_weight[0][78] , \input_weight[0][77] ,
         \input_weight[0][76] , \input_weight[0][75] , \input_weight[0][74] ,
         \input_weight[0][73] , \input_weight[0][72] , \input_weight[0][71] ,
         \input_weight[0][70] , \input_weight[0][69] , \input_weight[0][68] ,
         \input_weight[0][67] , \input_weight[0][66] , \input_weight[0][65] ,
         \input_weight[0][64] , \input_weight[0][63] , \input_weight[0][62] ,
         \input_weight[0][61] , \input_weight[0][60] , \input_weight[0][59] ,
         \input_weight[0][58] , \input_weight[0][57] , \input_weight[0][56] ,
         \input_weight[0][55] , \input_weight[0][54] , \input_weight[0][53] ,
         \input_weight[0][52] , \input_weight[0][51] , \input_weight[0][50] ,
         \input_weight[0][49] , \input_weight[0][48] , \input_weight[0][47] ,
         \input_weight[0][46] , \input_weight[0][45] , \input_weight[0][44] ,
         \input_weight[0][43] , \input_weight[0][42] , \input_weight[0][41] ,
         \input_weight[0][40] , \input_weight[0][39] , \input_weight[0][38] ,
         \input_weight[0][37] , \input_weight[0][36] , \input_weight[0][35] ,
         \input_weight[0][34] , \input_weight[0][33] , \input_weight[0][32] ,
         \input_weight[0][31] , \input_weight[0][30] , \input_weight[0][29] ,
         \input_weight[0][28] , \input_weight[0][27] , \input_weight[0][26] ,
         \input_weight[0][25] , \input_weight[0][24] , \input_weight[0][23] ,
         \input_weight[0][22] , \input_weight[0][21] , \input_weight[0][20] ,
         \input_weight[0][19] , \input_weight[0][18] , \input_weight[0][17] ,
         \input_weight[0][16] , \input_weight[0][15] , \input_weight[0][14] ,
         \input_weight[0][13] , \input_weight[0][12] , \input_weight[0][11] ,
         \input_weight[0][10] , \input_weight[0][9] , \input_weight[0][8] ,
         \input_weight[0][7] , \input_weight[0][6] , \input_weight[0][5] ,
         \input_weight[0][4] , \input_weight[0][3] , \input_weight[0][2] ,
         \input_weight[0][1] , \input_weight[0][0] , \input_bias[7][15] ,
         \input_bias[7][14] , \input_bias[7][13] , \input_bias[7][12] ,
         \input_bias[7][11] , \input_bias[7][10] , \input_bias[7][9] ,
         \input_bias[7][8] , \input_bias[7][7] , \input_bias[7][6] ,
         \input_bias[7][5] , \input_bias[7][4] , \input_bias[7][3] ,
         \input_bias[7][2] , \input_bias[7][1] , \input_bias[7][0] ,
         \input_bias[6][15] , \input_bias[6][14] , \input_bias[6][13] ,
         \input_bias[6][12] , \input_bias[6][11] , \input_bias[6][10] ,
         \input_bias[6][9] , \input_bias[6][8] , \input_bias[6][7] ,
         \input_bias[6][6] , \input_bias[6][5] , \input_bias[6][4] ,
         \input_bias[6][3] , \input_bias[6][2] , \input_bias[6][1] ,
         \input_bias[6][0] , \input_bias[5][15] , \input_bias[5][14] ,
         \input_bias[5][13] , \input_bias[5][12] , \input_bias[5][11] ,
         \input_bias[5][10] , \input_bias[5][9] , \input_bias[5][8] ,
         \input_bias[5][7] , \input_bias[5][6] , \input_bias[5][5] ,
         \input_bias[5][4] , \input_bias[5][3] , \input_bias[5][2] ,
         \input_bias[5][1] , \input_bias[5][0] , \input_bias[4][15] ,
         \input_bias[4][14] , \input_bias[4][13] , \input_bias[4][12] ,
         \input_bias[4][11] , \input_bias[4][10] , \input_bias[4][9] ,
         \input_bias[4][8] , \input_bias[4][7] , \input_bias[4][6] ,
         \input_bias[4][5] , \input_bias[4][4] , \input_bias[4][3] ,
         \input_bias[4][2] , \input_bias[4][1] , \input_bias[4][0] ,
         \input_bias[3][15] , \input_bias[3][14] , \input_bias[3][13] ,
         \input_bias[3][12] , \input_bias[3][11] , \input_bias[3][10] ,
         \input_bias[3][9] , \input_bias[3][8] , \input_bias[3][7] ,
         \input_bias[3][6] , \input_bias[3][5] , \input_bias[3][4] ,
         \input_bias[3][3] , \input_bias[3][2] , \input_bias[3][1] ,
         \input_bias[3][0] , \input_bias[2][15] , \input_bias[2][14] ,
         \input_bias[2][13] , \input_bias[2][12] , \input_bias[2][11] ,
         \input_bias[2][10] , \input_bias[2][9] , \input_bias[2][8] ,
         \input_bias[2][7] , \input_bias[2][6] , \input_bias[2][5] ,
         \input_bias[2][4] , \input_bias[2][3] , \input_bias[2][2] ,
         \input_bias[2][1] , \input_bias[2][0] , \input_bias[1][15] ,
         \input_bias[1][14] , \input_bias[1][13] , \input_bias[1][12] ,
         \input_bias[1][11] , \input_bias[1][10] , \input_bias[1][9] ,
         \input_bias[1][8] , \input_bias[1][7] , \input_bias[1][6] ,
         \input_bias[1][5] , \input_bias[1][4] , \input_bias[1][3] ,
         \input_bias[1][2] , \input_bias[1][1] , \input_bias[1][0] ,
         \input_bias[0][15] , \input_bias[0][14] , \input_bias[0][13] ,
         \input_bias[0][12] , \input_bias[0][11] , \input_bias[0][10] ,
         \input_bias[0][9] , \input_bias[0][8] , \input_bias[0][7] ,
         \input_bias[0][6] , \input_bias[0][5] , \input_bias[0][4] ,
         \input_bias[0][3] , \input_bias[0][2] , \input_bias[0][1] ,
         \input_bias[0][0] , N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N156, N312, N313, N314, N315, N317, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N428, N430, N432,
         N434, N436, N438, N440, N442, N444, N446, N448, N450, N452, N454,
         N456, N458, N460, N477, N478, N479, N480, N481, N482, N483, N484,
         \U3/U1/Z_5 , n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585;
  wire   [3:0] cur_state;
  wire   [15:0] neuron_BAR;
  wire   [3:0] nxt_state;
  wire   [3:0] mem_cur_state;
  wire   [3:0] mem_nxt_state;
  tri   [159:0] layer_data_out;
  tri   rst;
  tri   [7:0] done;
  tri   \output_value[7][15] ;
  tri   \output_value[7][14] ;
  tri   \output_value[7][13] ;
  tri   \output_value[7][12] ;
  tri   \output_value[7][11] ;
  tri   \output_value[7][10] ;
  tri   \output_value[7][9] ;
  tri   \output_value[7][8] ;
  tri   \output_value[7][7] ;
  tri   \output_value[7][6] ;
  tri   \output_value[7][5] ;
  tri   \output_value[7][4] ;
  tri   \output_value[7][3] ;
  tri   \output_value[7][2] ;
  tri   \output_value[7][1] ;
  tri   \output_value[7][0] ;
  tri   \output_value[6][15] ;
  tri   \output_value[6][14] ;
  tri   \output_value[6][13] ;
  tri   \output_value[6][12] ;
  tri   \output_value[6][11] ;
  tri   \output_value[6][10] ;
  tri   \output_value[6][9] ;
  tri   \output_value[6][8] ;
  tri   \output_value[6][7] ;
  tri   \output_value[6][6] ;
  tri   \output_value[6][5] ;
  tri   \output_value[6][4] ;
  tri   \output_value[6][3] ;
  tri   \output_value[6][2] ;
  tri   \output_value[6][1] ;
  tri   \output_value[6][0] ;
  tri   \output_value[5][15] ;
  tri   \output_value[5][14] ;
  tri   \output_value[5][13] ;
  tri   \output_value[5][12] ;
  tri   \output_value[5][11] ;
  tri   \output_value[5][10] ;
  tri   \output_value[5][9] ;
  tri   \output_value[5][8] ;
  tri   \output_value[5][7] ;
  tri   \output_value[5][6] ;
  tri   \output_value[5][5] ;
  tri   \output_value[5][4] ;
  tri   \output_value[5][3] ;
  tri   \output_value[5][2] ;
  tri   \output_value[5][1] ;
  tri   \output_value[5][0] ;
  tri   \output_value[4][15] ;
  tri   \output_value[4][14] ;
  tri   \output_value[4][13] ;
  tri   \output_value[4][12] ;
  tri   \output_value[4][11] ;
  tri   \output_value[4][10] ;
  tri   \output_value[4][9] ;
  tri   \output_value[4][8] ;
  tri   \output_value[4][7] ;
  tri   \output_value[4][6] ;
  tri   \output_value[4][5] ;
  tri   \output_value[4][4] ;
  tri   \output_value[4][3] ;
  tri   \output_value[4][2] ;
  tri   \output_value[4][1] ;
  tri   \output_value[4][0] ;
  tri   \output_value[3][15] ;
  tri   \output_value[3][14] ;
  tri   \output_value[3][13] ;
  tri   \output_value[3][12] ;
  tri   \output_value[3][11] ;
  tri   \output_value[3][10] ;
  tri   \output_value[3][9] ;
  tri   \output_value[3][8] ;
  tri   \output_value[3][7] ;
  tri   \output_value[3][6] ;
  tri   \output_value[3][5] ;
  tri   \output_value[3][4] ;
  tri   \output_value[3][3] ;
  tri   \output_value[3][2] ;
  tri   \output_value[3][1] ;
  tri   \output_value[3][0] ;
  tri   \output_value[2][15] ;
  tri   \output_value[2][14] ;
  tri   \output_value[2][13] ;
  tri   \output_value[2][12] ;
  tri   \output_value[2][11] ;
  tri   \output_value[2][10] ;
  tri   \output_value[2][9] ;
  tri   \output_value[2][8] ;
  tri   \output_value[2][7] ;
  tri   \output_value[2][6] ;
  tri   \output_value[2][5] ;
  tri   \output_value[2][4] ;
  tri   \output_value[2][3] ;
  tri   \output_value[2][2] ;
  tri   \output_value[2][1] ;
  tri   \output_value[2][0] ;
  tri   \output_value[1][15] ;
  tri   \output_value[1][14] ;
  tri   \output_value[1][13] ;
  tri   \output_value[1][12] ;
  tri   \output_value[1][11] ;
  tri   \output_value[1][10] ;
  tri   \output_value[1][9] ;
  tri   \output_value[1][8] ;
  tri   \output_value[1][7] ;
  tri   \output_value[1][6] ;
  tri   \output_value[1][5] ;
  tri   \output_value[1][4] ;
  tri   \output_value[1][3] ;
  tri   \output_value[1][2] ;
  tri   \output_value[1][1] ;
  tri   \output_value[1][0] ;
  tri   \output_value[0][15] ;
  tri   \output_value[0][14] ;
  tri   \output_value[0][13] ;
  tri   \output_value[0][12] ;
  tri   \output_value[0][11] ;
  tri   \output_value[0][10] ;
  tri   \output_value[0][9] ;
  tri   \output_value[0][8] ;
  tri   \output_value[0][7] ;
  tri   \output_value[0][6] ;
  tri   \output_value[0][5] ;
  tri   \output_value[0][4] ;
  tri   \output_value[0][3] ;
  tri   \output_value[0][2] ;
  tri   \output_value[0][1] ;
  tri   \output_value[0][0] ;
  tri   \forward_network[7][31] ;
  tri   \forward_network[7][30] ;
  tri   \forward_network[7][29] ;
  tri   \forward_network[7][28] ;
  tri   \forward_network[7][27] ;
  tri   \forward_network[7][26] ;
  tri   \forward_network[7][25] ;
  tri   \forward_network[7][24] ;
  tri   \forward_network[7][23] ;
  tri   \forward_network[7][22] ;
  tri   \forward_network[7][21] ;
  tri   \forward_network[7][20] ;
  tri   \forward_network[7][19] ;
  tri   \forward_network[7][18] ;
  tri   \forward_network[7][17] ;
  tri   \forward_network[7][16] ;
  tri   \forward_network[7][15] ;
  tri   \forward_network[7][14] ;
  tri   \forward_network[7][13] ;
  tri   \forward_network[7][12] ;
  tri   \forward_network[7][11] ;
  tri   \forward_network[7][10] ;
  tri   \forward_network[7][9] ;
  tri   \forward_network[7][8] ;
  tri   \forward_network[7][7] ;
  tri   \forward_network[7][6] ;
  tri   \forward_network[7][5] ;
  tri   \forward_network[7][4] ;
  tri   \forward_network[7][3] ;
  tri   \forward_network[7][2] ;
  tri   \forward_network[7][1] ;
  tri   \forward_network[7][0] ;
  tri   \forward_network[6][31] ;
  tri   \forward_network[6][30] ;
  tri   \forward_network[6][29] ;
  tri   \forward_network[6][28] ;
  tri   \forward_network[6][27] ;
  tri   \forward_network[6][26] ;
  tri   \forward_network[6][25] ;
  tri   \forward_network[6][24] ;
  tri   \forward_network[6][23] ;
  tri   \forward_network[6][22] ;
  tri   \forward_network[6][21] ;
  tri   \forward_network[6][20] ;
  tri   \forward_network[6][19] ;
  tri   \forward_network[6][18] ;
  tri   \forward_network[6][17] ;
  tri   \forward_network[6][16] ;
  tri   \forward_network[6][15] ;
  tri   \forward_network[6][14] ;
  tri   \forward_network[6][13] ;
  tri   \forward_network[6][12] ;
  tri   \forward_network[6][11] ;
  tri   \forward_network[6][10] ;
  tri   \forward_network[6][9] ;
  tri   \forward_network[6][8] ;
  tri   \forward_network[6][7] ;
  tri   \forward_network[6][6] ;
  tri   \forward_network[6][5] ;
  tri   \forward_network[6][4] ;
  tri   \forward_network[6][3] ;
  tri   \forward_network[6][2] ;
  tri   \forward_network[6][1] ;
  tri   \forward_network[6][0] ;
  tri   \forward_network[5][31] ;
  tri   \forward_network[5][30] ;
  tri   \forward_network[5][29] ;
  tri   \forward_network[5][28] ;
  tri   \forward_network[5][27] ;
  tri   \forward_network[5][26] ;
  tri   \forward_network[5][25] ;
  tri   \forward_network[5][24] ;
  tri   \forward_network[5][23] ;
  tri   \forward_network[5][22] ;
  tri   \forward_network[5][21] ;
  tri   \forward_network[5][20] ;
  tri   \forward_network[5][19] ;
  tri   \forward_network[5][18] ;
  tri   \forward_network[5][17] ;
  tri   \forward_network[5][16] ;
  tri   \forward_network[5][15] ;
  tri   \forward_network[5][14] ;
  tri   \forward_network[5][13] ;
  tri   \forward_network[5][12] ;
  tri   \forward_network[5][11] ;
  tri   \forward_network[5][10] ;
  tri   \forward_network[5][9] ;
  tri   \forward_network[5][8] ;
  tri   \forward_network[5][7] ;
  tri   \forward_network[5][6] ;
  tri   \forward_network[5][5] ;
  tri   \forward_network[5][4] ;
  tri   \forward_network[5][3] ;
  tri   \forward_network[5][2] ;
  tri   \forward_network[5][1] ;
  tri   \forward_network[5][0] ;
  tri   \forward_network[4][31] ;
  tri   \forward_network[4][30] ;
  tri   \forward_network[4][29] ;
  tri   \forward_network[4][28] ;
  tri   \forward_network[4][27] ;
  tri   \forward_network[4][26] ;
  tri   \forward_network[4][25] ;
  tri   \forward_network[4][24] ;
  tri   \forward_network[4][23] ;
  tri   \forward_network[4][22] ;
  tri   \forward_network[4][21] ;
  tri   \forward_network[4][20] ;
  tri   \forward_network[4][19] ;
  tri   \forward_network[4][18] ;
  tri   \forward_network[4][17] ;
  tri   \forward_network[4][16] ;
  tri   \forward_network[4][15] ;
  tri   \forward_network[4][14] ;
  tri   \forward_network[4][13] ;
  tri   \forward_network[4][12] ;
  tri   \forward_network[4][11] ;
  tri   \forward_network[4][10] ;
  tri   \forward_network[4][9] ;
  tri   \forward_network[4][8] ;
  tri   \forward_network[4][7] ;
  tri   \forward_network[4][6] ;
  tri   \forward_network[4][5] ;
  tri   \forward_network[4][4] ;
  tri   \forward_network[4][3] ;
  tri   \forward_network[4][2] ;
  tri   \forward_network[4][1] ;
  tri   \forward_network[4][0] ;
  tri   \forward_network[3][31] ;
  tri   \forward_network[3][30] ;
  tri   \forward_network[3][29] ;
  tri   \forward_network[3][28] ;
  tri   \forward_network[3][27] ;
  tri   \forward_network[3][26] ;
  tri   \forward_network[3][25] ;
  tri   \forward_network[3][24] ;
  tri   \forward_network[3][23] ;
  tri   \forward_network[3][22] ;
  tri   \forward_network[3][21] ;
  tri   \forward_network[3][20] ;
  tri   \forward_network[3][19] ;
  tri   \forward_network[3][18] ;
  tri   \forward_network[3][17] ;
  tri   \forward_network[3][16] ;
  tri   \forward_network[3][15] ;
  tri   \forward_network[3][14] ;
  tri   \forward_network[3][13] ;
  tri   \forward_network[3][12] ;
  tri   \forward_network[3][11] ;
  tri   \forward_network[3][10] ;
  tri   \forward_network[3][9] ;
  tri   \forward_network[3][8] ;
  tri   \forward_network[3][7] ;
  tri   \forward_network[3][6] ;
  tri   \forward_network[3][5] ;
  tri   \forward_network[3][4] ;
  tri   \forward_network[3][3] ;
  tri   \forward_network[3][2] ;
  tri   \forward_network[3][1] ;
  tri   \forward_network[3][0] ;
  tri   \forward_network[2][31] ;
  tri   \forward_network[2][30] ;
  tri   \forward_network[2][29] ;
  tri   \forward_network[2][28] ;
  tri   \forward_network[2][27] ;
  tri   \forward_network[2][26] ;
  tri   \forward_network[2][25] ;
  tri   \forward_network[2][24] ;
  tri   \forward_network[2][23] ;
  tri   \forward_network[2][22] ;
  tri   \forward_network[2][21] ;
  tri   \forward_network[2][20] ;
  tri   \forward_network[2][19] ;
  tri   \forward_network[2][18] ;
  tri   \forward_network[2][17] ;
  tri   \forward_network[2][16] ;
  tri   \forward_network[2][15] ;
  tri   \forward_network[2][14] ;
  tri   \forward_network[2][13] ;
  tri   \forward_network[2][12] ;
  tri   \forward_network[2][11] ;
  tri   \forward_network[2][10] ;
  tri   \forward_network[2][9] ;
  tri   \forward_network[2][8] ;
  tri   \forward_network[2][7] ;
  tri   \forward_network[2][6] ;
  tri   \forward_network[2][5] ;
  tri   \forward_network[2][4] ;
  tri   \forward_network[2][3] ;
  tri   \forward_network[2][2] ;
  tri   \forward_network[2][1] ;
  tri   \forward_network[2][0] ;
  tri   \forward_network[1][31] ;
  tri   \forward_network[1][30] ;
  tri   \forward_network[1][29] ;
  tri   \forward_network[1][28] ;
  tri   \forward_network[1][27] ;
  tri   \forward_network[1][26] ;
  tri   \forward_network[1][25] ;
  tri   \forward_network[1][24] ;
  tri   \forward_network[1][23] ;
  tri   \forward_network[1][22] ;
  tri   \forward_network[1][21] ;
  tri   \forward_network[1][20] ;
  tri   \forward_network[1][19] ;
  tri   \forward_network[1][18] ;
  tri   \forward_network[1][17] ;
  tri   \forward_network[1][16] ;
  tri   \forward_network[1][15] ;
  tri   \forward_network[1][14] ;
  tri   \forward_network[1][13] ;
  tri   \forward_network[1][12] ;
  tri   \forward_network[1][11] ;
  tri   \forward_network[1][10] ;
  tri   \forward_network[1][9] ;
  tri   \forward_network[1][8] ;
  tri   \forward_network[1][7] ;
  tri   \forward_network[1][6] ;
  tri   \forward_network[1][5] ;
  tri   \forward_network[1][4] ;
  tri   \forward_network[1][3] ;
  tri   \forward_network[1][2] ;
  tri   \forward_network[1][1] ;
  tri   \forward_network[1][0] ;
  tri   \forward_network[0][31] ;
  tri   \forward_network[0][30] ;
  tri   \forward_network[0][29] ;
  tri   \forward_network[0][28] ;
  tri   \forward_network[0][27] ;
  tri   \forward_network[0][26] ;
  tri   \forward_network[0][25] ;
  tri   \forward_network[0][24] ;
  tri   \forward_network[0][23] ;
  tri   \forward_network[0][22] ;
  tri   \forward_network[0][21] ;
  tri   \forward_network[0][20] ;
  tri   \forward_network[0][19] ;
  tri   \forward_network[0][18] ;
  tri   \forward_network[0][17] ;
  tri   \forward_network[0][16] ;
  tri   \forward_network[0][15] ;
  tri   \forward_network[0][14] ;
  tri   \forward_network[0][13] ;
  tri   \forward_network[0][12] ;
  tri   \forward_network[0][11] ;
  tri   \forward_network[0][10] ;
  tri   \forward_network[0][9] ;
  tri   \forward_network[0][8] ;
  tri   \forward_network[0][7] ;
  tri   \forward_network[0][6] ;
  tri   \forward_network[0][5] ;
  tri   \forward_network[0][4] ;
  tri   \forward_network[0][3] ;
  tri   \forward_network[0][2] ;
  tri   \forward_network[0][1] ;
  tri   \forward_network[0][0] ;
  tri   [19:0] fwd_routing_engine_control;
  tri   fwd_routing_engine_done;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;
  assign layer_done = RE;

  EDFQD2 \len_reg[0]  ( .D(n584), .E(N312), .CP(clk), .Q(len[0]) );
  EDFQD2 \len_reg[1]  ( .D(N313), .E(N312), .CP(clk), .Q(len[1]) );
  EDFQD2 \len_reg[2]  ( .D(N313), .E(N312), .CP(clk), .Q(len[2]) );
  EDFQD2 \len_reg[3]  ( .D(N313), .E(N312), .CP(clk), .Q(len[3]) );
  EDFQD2 \addr_reg[0]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[0]) );
  EDFQD2 \addr_reg[1]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[1]) );
  EDFQD2 \addr_reg[2]  ( .D(N320), .E(N312), .CP(clk), .Q(addr[2]) );
  EDFQD2 \addr_reg[3]  ( .D(N321), .E(N312), .CP(clk), .Q(addr[3]) );
  EDFQD2 \addr_reg[4]  ( .D(N322), .E(N312), .CP(clk), .Q(addr[4]) );
  EDFQD2 \addr_reg[5]  ( .D(N323), .E(N312), .CP(clk), .Q(addr[5]) );
  EDFQD2 \addr_reg[6]  ( .D(N324), .E(N312), .CP(clk), .Q(addr[6]) );
  EDFQD2 \addr_reg[7]  ( .D(N325), .E(N312), .CP(clk), .Q(addr[7]) );
  EDFQD2 \addr_reg[8]  ( .D(N326), .E(N312), .CP(clk), .Q(addr[8]) );
  EDFQD2 \addr_reg[9]  ( .D(N327), .E(N312), .CP(clk), .Q(addr[9]) );
  EDFQD2 \addr_reg[10]  ( .D(N328), .E(N312), .CP(clk), .Q(addr[10]) );
  EDFQD2 \addr_reg[11]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[11]) );
  EDFQD2 \addr_reg[12]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[12]) );
  EDFQD2 \addr_reg[13]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[13]) );
  EDFQD2 \addr_reg[14]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[14]) );
  EDFQD2 \addr_reg[15]  ( .D(WE), .E(N312), .CP(clk), .Q(addr[15]) );
  neuron_0 \generate_neurons[0].u_neuron  ( .input_value({
        \input_value[0][127] , \input_value[0][126] , \input_value[0][125] , 
        \input_value[0][124] , \input_value[0][123] , \input_value[0][122] , 
        \input_value[0][121] , \input_value[0][120] , \input_value[0][119] , 
        \input_value[0][118] , \input_value[0][117] , \input_value[0][116] , 
        \input_value[0][115] , \input_value[0][114] , \input_value[0][113] , 
        \input_value[0][112] , \input_value[0][111] , \input_value[0][110] , 
        \input_value[0][109] , \input_value[0][108] , \input_value[0][107] , 
        \input_value[0][106] , \input_value[0][105] , \input_value[0][104] , 
        \input_value[0][103] , \input_value[0][102] , \input_value[0][101] , 
        \input_value[0][100] , \input_value[0][99] , \input_value[0][98] , 
        \input_value[0][97] , \input_value[0][96] , \input_value[0][95] , 
        \input_value[0][94] , \input_value[0][93] , \input_value[0][92] , 
        \input_value[0][91] , \input_value[0][90] , \input_value[0][89] , 
        \input_value[0][88] , \input_value[0][87] , \input_value[0][86] , 
        \input_value[0][85] , \input_value[0][84] , \input_value[0][83] , 
        \input_value[0][82] , \input_value[0][81] , \input_value[0][80] , 
        \input_value[0][79] , \input_value[0][78] , \input_value[0][77] , 
        \input_value[0][76] , \input_value[0][75] , \input_value[0][74] , 
        \input_value[0][73] , \input_value[0][72] , \input_value[0][71] , 
        \input_value[0][70] , \input_value[0][69] , \input_value[0][68] , 
        \input_value[0][67] , \input_value[0][66] , \input_value[0][65] , 
        \input_value[0][64] , \input_value[0][63] , \input_value[0][62] , 
        \input_value[0][61] , \input_value[0][60] , \input_value[0][59] , 
        \input_value[0][58] , \input_value[0][57] , \input_value[0][56] , 
        \input_value[0][55] , \input_value[0][54] , \input_value[0][53] , 
        \input_value[0][52] , \input_value[0][51] , \input_value[0][50] , 
        \input_value[0][49] , \input_value[0][48] , \input_value[0][47] , 
        \input_value[0][46] , \input_value[0][45] , \input_value[0][44] , 
        \input_value[0][43] , \input_value[0][42] , \input_value[0][41] , 
        \input_value[0][40] , \input_value[0][39] , \input_value[0][38] , 
        \input_value[0][37] , \input_value[0][36] , \input_value[0][35] , 
        \input_value[0][34] , \input_value[0][33] , \input_value[0][32] , 
        \input_value[0][31] , \input_value[0][30] , \input_value[0][29] , 
        \input_value[0][28] , \input_value[0][27] , \input_value[0][26] , 
        \input_value[0][25] , \input_value[0][24] , \input_value[0][23] , 
        \input_value[0][22] , \input_value[0][21] , \input_value[0][20] , 
        \input_value[0][19] , \input_value[0][18] , \input_value[0][17] , 
        \input_value[0][16] , \input_value[0][15] , \input_value[0][14] , 
        \input_value[0][13] , \input_value[0][12] , \input_value[0][11] , 
        \input_value[0][10] , \input_value[0][9] , \input_value[0][8] , 
        \input_value[0][7] , \input_value[0][6] , \input_value[0][5] , 
        \input_value[0][4] , \input_value[0][3] , \input_value[0][2] , 
        \input_value[0][1] , \input_value[0][0] }), .input_weight({
        \input_weight[0][127] , \input_weight[0][126] , \input_weight[0][125] , 
        \input_weight[0][124] , \input_weight[0][123] , \input_weight[0][122] , 
        \input_weight[0][121] , \input_weight[0][120] , \input_weight[0][119] , 
        \input_weight[0][118] , \input_weight[0][117] , \input_weight[0][116] , 
        \input_weight[0][115] , \input_weight[0][114] , \input_weight[0][113] , 
        \input_weight[0][112] , \input_weight[0][111] , \input_weight[0][110] , 
        \input_weight[0][109] , \input_weight[0][108] , \input_weight[0][107] , 
        \input_weight[0][106] , \input_weight[0][105] , \input_weight[0][104] , 
        \input_weight[0][103] , \input_weight[0][102] , \input_weight[0][101] , 
        \input_weight[0][100] , \input_weight[0][99] , \input_weight[0][98] , 
        \input_weight[0][97] , \input_weight[0][96] , \input_weight[0][95] , 
        \input_weight[0][94] , \input_weight[0][93] , \input_weight[0][92] , 
        \input_weight[0][91] , \input_weight[0][90] , \input_weight[0][89] , 
        \input_weight[0][88] , \input_weight[0][87] , \input_weight[0][86] , 
        \input_weight[0][85] , \input_weight[0][84] , \input_weight[0][83] , 
        \input_weight[0][82] , \input_weight[0][81] , \input_weight[0][80] , 
        \input_weight[0][79] , \input_weight[0][78] , \input_weight[0][77] , 
        \input_weight[0][76] , \input_weight[0][75] , \input_weight[0][74] , 
        \input_weight[0][73] , \input_weight[0][72] , \input_weight[0][71] , 
        \input_weight[0][70] , \input_weight[0][69] , \input_weight[0][68] , 
        \input_weight[0][67] , \input_weight[0][66] , \input_weight[0][65] , 
        \input_weight[0][64] , \input_weight[0][63] , \input_weight[0][62] , 
        \input_weight[0][61] , \input_weight[0][60] , \input_weight[0][59] , 
        \input_weight[0][58] , \input_weight[0][57] , \input_weight[0][56] , 
        \input_weight[0][55] , \input_weight[0][54] , \input_weight[0][53] , 
        \input_weight[0][52] , \input_weight[0][51] , \input_weight[0][50] , 
        \input_weight[0][49] , \input_weight[0][48] , \input_weight[0][47] , 
        \input_weight[0][46] , \input_weight[0][45] , \input_weight[0][44] , 
        \input_weight[0][43] , \input_weight[0][42] , \input_weight[0][41] , 
        \input_weight[0][40] , \input_weight[0][39] , \input_weight[0][38] , 
        \input_weight[0][37] , \input_weight[0][36] , \input_weight[0][35] , 
        \input_weight[0][34] , \input_weight[0][33] , \input_weight[0][32] , 
        \input_weight[0][31] , \input_weight[0][30] , \input_weight[0][29] , 
        \input_weight[0][28] , \input_weight[0][27] , \input_weight[0][26] , 
        \input_weight[0][25] , \input_weight[0][24] , \input_weight[0][23] , 
        \input_weight[0][22] , \input_weight[0][21] , \input_weight[0][20] , 
        \input_weight[0][19] , \input_weight[0][18] , \input_weight[0][17] , 
        \input_weight[0][16] , \input_weight[0][15] , \input_weight[0][14] , 
        \input_weight[0][13] , \input_weight[0][12] , \input_weight[0][11] , 
        \input_weight[0][10] , \input_weight[0][9] , \input_weight[0][8] , 
        \input_weight[0][7] , \input_weight[0][6] , \input_weight[0][5] , 
        \input_weight[0][4] , \input_weight[0][3] , \input_weight[0][2] , 
        \input_weight[0][1] , \input_weight[0][0] }), .input_bias({
        \input_bias[0][15] , \input_bias[0][14] , \input_bias[0][13] , 
        \input_bias[0][12] , \input_bias[0][11] , \input_bias[0][10] , 
        \input_bias[0][9] , \input_bias[0][8] , \input_bias[0][7] , 
        \input_bias[0][6] , \input_bias[0][5] , \input_bias[0][4] , 
        \input_bias[0][3] , \input_bias[0][2] , \input_bias[0][1] , 
        \input_bias[0][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[0][15] , \output_value[0][14] , \output_value[0][13] , 
        \output_value[0][12] , \output_value[0][11] , \output_value[0][10] , 
        \output_value[0][9] , \output_value[0][8] , \output_value[0][7] , 
        \output_value[0][6] , \output_value[0][5] , \output_value[0][4] , 
        \output_value[0][3] , \output_value[0][2] , \output_value[0][1] , 
        \output_value[0][0] }), .clk(WE) );
  neuron_7 \generate_neurons[1].u_neuron  ( .input_value({
        \input_value[1][127] , \input_value[1][126] , \input_value[1][125] , 
        \input_value[1][124] , \input_value[1][123] , \input_value[1][122] , 
        \input_value[1][121] , \input_value[1][120] , \input_value[1][119] , 
        \input_value[1][118] , \input_value[1][117] , \input_value[1][116] , 
        \input_value[1][115] , \input_value[1][114] , \input_value[1][113] , 
        \input_value[1][112] , \input_value[1][111] , \input_value[1][110] , 
        \input_value[1][109] , \input_value[1][108] , \input_value[1][107] , 
        \input_value[1][106] , \input_value[1][105] , \input_value[1][104] , 
        \input_value[1][103] , \input_value[1][102] , \input_value[1][101] , 
        \input_value[1][100] , \input_value[1][99] , \input_value[1][98] , 
        \input_value[1][97] , \input_value[1][96] , \input_value[1][95] , 
        \input_value[1][94] , \input_value[1][93] , \input_value[1][92] , 
        \input_value[1][91] , \input_value[1][90] , \input_value[1][89] , 
        \input_value[1][88] , \input_value[1][87] , \input_value[1][86] , 
        \input_value[1][85] , \input_value[1][84] , \input_value[1][83] , 
        \input_value[1][82] , \input_value[1][81] , \input_value[1][80] , 
        \input_value[1][79] , \input_value[1][78] , \input_value[1][77] , 
        \input_value[1][76] , \input_value[1][75] , \input_value[1][74] , 
        \input_value[1][73] , \input_value[1][72] , \input_value[1][71] , 
        \input_value[1][70] , \input_value[1][69] , \input_value[1][68] , 
        \input_value[1][67] , \input_value[1][66] , \input_value[1][65] , 
        \input_value[1][64] , \input_value[1][63] , \input_value[1][62] , 
        \input_value[1][61] , \input_value[1][60] , \input_value[1][59] , 
        \input_value[1][58] , \input_value[1][57] , \input_value[1][56] , 
        \input_value[1][55] , \input_value[1][54] , \input_value[1][53] , 
        \input_value[1][52] , \input_value[1][51] , \input_value[1][50] , 
        \input_value[1][49] , \input_value[1][48] , \input_value[1][47] , 
        \input_value[1][46] , \input_value[1][45] , \input_value[1][44] , 
        \input_value[1][43] , \input_value[1][42] , \input_value[1][41] , 
        \input_value[1][40] , \input_value[1][39] , \input_value[1][38] , 
        \input_value[1][37] , \input_value[1][36] , \input_value[1][35] , 
        \input_value[1][34] , \input_value[1][33] , \input_value[1][32] , 
        \input_value[1][31] , \input_value[1][30] , \input_value[1][29] , 
        \input_value[1][28] , \input_value[1][27] , \input_value[1][26] , 
        \input_value[1][25] , \input_value[1][24] , \input_value[1][23] , 
        \input_value[1][22] , \input_value[1][21] , \input_value[1][20] , 
        \input_value[1][19] , \input_value[1][18] , \input_value[1][17] , 
        \input_value[1][16] , \input_value[1][15] , \input_value[1][14] , 
        \input_value[1][13] , \input_value[1][12] , \input_value[1][11] , 
        \input_value[1][10] , \input_value[1][9] , \input_value[1][8] , 
        \input_value[1][7] , \input_value[1][6] , \input_value[1][5] , 
        \input_value[1][4] , \input_value[1][3] , \input_value[1][2] , 
        \input_value[1][1] , \input_value[1][0] }), .input_weight({
        \input_weight[1][127] , \input_weight[1][126] , \input_weight[1][125] , 
        \input_weight[1][124] , \input_weight[1][123] , \input_weight[1][122] , 
        \input_weight[1][121] , \input_weight[1][120] , \input_weight[1][119] , 
        \input_weight[1][118] , \input_weight[1][117] , \input_weight[1][116] , 
        \input_weight[1][115] , \input_weight[1][114] , \input_weight[1][113] , 
        \input_weight[1][112] , \input_weight[1][111] , \input_weight[1][110] , 
        \input_weight[1][109] , \input_weight[1][108] , \input_weight[1][107] , 
        \input_weight[1][106] , \input_weight[1][105] , \input_weight[1][104] , 
        \input_weight[1][103] , \input_weight[1][102] , \input_weight[1][101] , 
        \input_weight[1][100] , \input_weight[1][99] , \input_weight[1][98] , 
        \input_weight[1][97] , \input_weight[1][96] , \input_weight[1][95] , 
        \input_weight[1][94] , \input_weight[1][93] , \input_weight[1][92] , 
        \input_weight[1][91] , \input_weight[1][90] , \input_weight[1][89] , 
        \input_weight[1][88] , \input_weight[1][87] , \input_weight[1][86] , 
        \input_weight[1][85] , \input_weight[1][84] , \input_weight[1][83] , 
        \input_weight[1][82] , \input_weight[1][81] , \input_weight[1][80] , 
        \input_weight[1][79] , \input_weight[1][78] , \input_weight[1][77] , 
        \input_weight[1][76] , \input_weight[1][75] , \input_weight[1][74] , 
        \input_weight[1][73] , \input_weight[1][72] , \input_weight[1][71] , 
        \input_weight[1][70] , \input_weight[1][69] , \input_weight[1][68] , 
        \input_weight[1][67] , \input_weight[1][66] , \input_weight[1][65] , 
        \input_weight[1][64] , \input_weight[1][63] , \input_weight[1][62] , 
        \input_weight[1][61] , \input_weight[1][60] , \input_weight[1][59] , 
        \input_weight[1][58] , \input_weight[1][57] , \input_weight[1][56] , 
        \input_weight[1][55] , \input_weight[1][54] , \input_weight[1][53] , 
        \input_weight[1][52] , \input_weight[1][51] , \input_weight[1][50] , 
        \input_weight[1][49] , \input_weight[1][48] , \input_weight[1][47] , 
        \input_weight[1][46] , \input_weight[1][45] , \input_weight[1][44] , 
        \input_weight[1][43] , \input_weight[1][42] , \input_weight[1][41] , 
        \input_weight[1][40] , \input_weight[1][39] , \input_weight[1][38] , 
        \input_weight[1][37] , \input_weight[1][36] , \input_weight[1][35] , 
        \input_weight[1][34] , \input_weight[1][33] , \input_weight[1][32] , 
        \input_weight[1][31] , \input_weight[1][30] , \input_weight[1][29] , 
        \input_weight[1][28] , \input_weight[1][27] , \input_weight[1][26] , 
        \input_weight[1][25] , \input_weight[1][24] , \input_weight[1][23] , 
        \input_weight[1][22] , \input_weight[1][21] , \input_weight[1][20] , 
        \input_weight[1][19] , \input_weight[1][18] , \input_weight[1][17] , 
        \input_weight[1][16] , \input_weight[1][15] , \input_weight[1][14] , 
        \input_weight[1][13] , \input_weight[1][12] , \input_weight[1][11] , 
        \input_weight[1][10] , \input_weight[1][9] , \input_weight[1][8] , 
        \input_weight[1][7] , \input_weight[1][6] , \input_weight[1][5] , 
        \input_weight[1][4] , \input_weight[1][3] , \input_weight[1][2] , 
        \input_weight[1][1] , \input_weight[1][0] }), .input_bias({
        \input_bias[1][15] , \input_bias[1][14] , \input_bias[1][13] , 
        \input_bias[1][12] , \input_bias[1][11] , \input_bias[1][10] , 
        \input_bias[1][9] , \input_bias[1][8] , \input_bias[1][7] , 
        \input_bias[1][6] , \input_bias[1][5] , \input_bias[1][4] , 
        \input_bias[1][3] , \input_bias[1][2] , \input_bias[1][1] , 
        \input_bias[1][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[1][15] , \output_value[1][14] , \output_value[1][13] , 
        \output_value[1][12] , \output_value[1][11] , \output_value[1][10] , 
        \output_value[1][9] , \output_value[1][8] , \output_value[1][7] , 
        \output_value[1][6] , \output_value[1][5] , \output_value[1][4] , 
        \output_value[1][3] , \output_value[1][2] , \output_value[1][1] , 
        \output_value[1][0] }), .clk(WE) );
  neuron_6 \generate_neurons[2].u_neuron  ( .input_value({
        \input_value[2][127] , \input_value[2][126] , \input_value[2][125] , 
        \input_value[2][124] , \input_value[2][123] , \input_value[2][122] , 
        \input_value[2][121] , \input_value[2][120] , \input_value[2][119] , 
        \input_value[2][118] , \input_value[2][117] , \input_value[2][116] , 
        \input_value[2][115] , \input_value[2][114] , \input_value[2][113] , 
        \input_value[2][112] , \input_value[2][111] , \input_value[2][110] , 
        \input_value[2][109] , \input_value[2][108] , \input_value[2][107] , 
        \input_value[2][106] , \input_value[2][105] , \input_value[2][104] , 
        \input_value[2][103] , \input_value[2][102] , \input_value[2][101] , 
        \input_value[2][100] , \input_value[2][99] , \input_value[2][98] , 
        \input_value[2][97] , \input_value[2][96] , \input_value[2][95] , 
        \input_value[2][94] , \input_value[2][93] , \input_value[2][92] , 
        \input_value[2][91] , \input_value[2][90] , \input_value[2][89] , 
        \input_value[2][88] , \input_value[2][87] , \input_value[2][86] , 
        \input_value[2][85] , \input_value[2][84] , \input_value[2][83] , 
        \input_value[2][82] , \input_value[2][81] , \input_value[2][80] , 
        \input_value[2][79] , \input_value[2][78] , \input_value[2][77] , 
        \input_value[2][76] , \input_value[2][75] , \input_value[2][74] , 
        \input_value[2][73] , \input_value[2][72] , \input_value[2][71] , 
        \input_value[2][70] , \input_value[2][69] , \input_value[2][68] , 
        \input_value[2][67] , \input_value[2][66] , \input_value[2][65] , 
        \input_value[2][64] , \input_value[2][63] , \input_value[2][62] , 
        \input_value[2][61] , \input_value[2][60] , \input_value[2][59] , 
        \input_value[2][58] , \input_value[2][57] , \input_value[2][56] , 
        \input_value[2][55] , \input_value[2][54] , \input_value[2][53] , 
        \input_value[2][52] , \input_value[2][51] , \input_value[2][50] , 
        \input_value[2][49] , \input_value[2][48] , \input_value[2][47] , 
        \input_value[2][46] , \input_value[2][45] , \input_value[2][44] , 
        \input_value[2][43] , \input_value[2][42] , \input_value[2][41] , 
        \input_value[2][40] , \input_value[2][39] , \input_value[2][38] , 
        \input_value[2][37] , \input_value[2][36] , \input_value[2][35] , 
        \input_value[2][34] , \input_value[2][33] , \input_value[2][32] , 
        \input_value[2][31] , \input_value[2][30] , \input_value[2][29] , 
        \input_value[2][28] , \input_value[2][27] , \input_value[2][26] , 
        \input_value[2][25] , \input_value[2][24] , \input_value[2][23] , 
        \input_value[2][22] , \input_value[2][21] , \input_value[2][20] , 
        \input_value[2][19] , \input_value[2][18] , \input_value[2][17] , 
        \input_value[2][16] , \input_value[2][15] , \input_value[2][14] , 
        \input_value[2][13] , \input_value[2][12] , \input_value[2][11] , 
        \input_value[2][10] , \input_value[2][9] , \input_value[2][8] , 
        \input_value[2][7] , \input_value[2][6] , \input_value[2][5] , 
        \input_value[2][4] , \input_value[2][3] , \input_value[2][2] , 
        \input_value[2][1] , \input_value[2][0] }), .input_weight({
        \input_weight[2][127] , \input_weight[2][126] , \input_weight[2][125] , 
        \input_weight[2][124] , \input_weight[2][123] , \input_weight[2][122] , 
        \input_weight[2][121] , \input_weight[2][120] , \input_weight[2][119] , 
        \input_weight[2][118] , \input_weight[2][117] , \input_weight[2][116] , 
        \input_weight[2][115] , \input_weight[2][114] , \input_weight[2][113] , 
        \input_weight[2][112] , \input_weight[2][111] , \input_weight[2][110] , 
        \input_weight[2][109] , \input_weight[2][108] , \input_weight[2][107] , 
        \input_weight[2][106] , \input_weight[2][105] , \input_weight[2][104] , 
        \input_weight[2][103] , \input_weight[2][102] , \input_weight[2][101] , 
        \input_weight[2][100] , \input_weight[2][99] , \input_weight[2][98] , 
        \input_weight[2][97] , \input_weight[2][96] , \input_weight[2][95] , 
        \input_weight[2][94] , \input_weight[2][93] , \input_weight[2][92] , 
        \input_weight[2][91] , \input_weight[2][90] , \input_weight[2][89] , 
        \input_weight[2][88] , \input_weight[2][87] , \input_weight[2][86] , 
        \input_weight[2][85] , \input_weight[2][84] , \input_weight[2][83] , 
        \input_weight[2][82] , \input_weight[2][81] , \input_weight[2][80] , 
        \input_weight[2][79] , \input_weight[2][78] , \input_weight[2][77] , 
        \input_weight[2][76] , \input_weight[2][75] , \input_weight[2][74] , 
        \input_weight[2][73] , \input_weight[2][72] , \input_weight[2][71] , 
        \input_weight[2][70] , \input_weight[2][69] , \input_weight[2][68] , 
        \input_weight[2][67] , \input_weight[2][66] , \input_weight[2][65] , 
        \input_weight[2][64] , \input_weight[2][63] , \input_weight[2][62] , 
        \input_weight[2][61] , \input_weight[2][60] , \input_weight[2][59] , 
        \input_weight[2][58] , \input_weight[2][57] , \input_weight[2][56] , 
        \input_weight[2][55] , \input_weight[2][54] , \input_weight[2][53] , 
        \input_weight[2][52] , \input_weight[2][51] , \input_weight[2][50] , 
        \input_weight[2][49] , \input_weight[2][48] , \input_weight[2][47] , 
        \input_weight[2][46] , \input_weight[2][45] , \input_weight[2][44] , 
        \input_weight[2][43] , \input_weight[2][42] , \input_weight[2][41] , 
        \input_weight[2][40] , \input_weight[2][39] , \input_weight[2][38] , 
        \input_weight[2][37] , \input_weight[2][36] , \input_weight[2][35] , 
        \input_weight[2][34] , \input_weight[2][33] , \input_weight[2][32] , 
        \input_weight[2][31] , \input_weight[2][30] , \input_weight[2][29] , 
        \input_weight[2][28] , \input_weight[2][27] , \input_weight[2][26] , 
        \input_weight[2][25] , \input_weight[2][24] , \input_weight[2][23] , 
        \input_weight[2][22] , \input_weight[2][21] , \input_weight[2][20] , 
        \input_weight[2][19] , \input_weight[2][18] , \input_weight[2][17] , 
        \input_weight[2][16] , \input_weight[2][15] , \input_weight[2][14] , 
        \input_weight[2][13] , \input_weight[2][12] , \input_weight[2][11] , 
        \input_weight[2][10] , \input_weight[2][9] , \input_weight[2][8] , 
        \input_weight[2][7] , \input_weight[2][6] , \input_weight[2][5] , 
        \input_weight[2][4] , \input_weight[2][3] , \input_weight[2][2] , 
        \input_weight[2][1] , \input_weight[2][0] }), .input_bias({
        \input_bias[2][15] , \input_bias[2][14] , \input_bias[2][13] , 
        \input_bias[2][12] , \input_bias[2][11] , \input_bias[2][10] , 
        \input_bias[2][9] , \input_bias[2][8] , \input_bias[2][7] , 
        \input_bias[2][6] , \input_bias[2][5] , \input_bias[2][4] , 
        \input_bias[2][3] , \input_bias[2][2] , \input_bias[2][1] , 
        \input_bias[2][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[2][15] , \output_value[2][14] , \output_value[2][13] , 
        \output_value[2][12] , \output_value[2][11] , \output_value[2][10] , 
        \output_value[2][9] , \output_value[2][8] , \output_value[2][7] , 
        \output_value[2][6] , \output_value[2][5] , \output_value[2][4] , 
        \output_value[2][3] , \output_value[2][2] , \output_value[2][1] , 
        \output_value[2][0] }), .clk(WE) );
  neuron_5 \generate_neurons[3].u_neuron  ( .input_value({
        \input_value[3][127] , \input_value[3][126] , \input_value[3][125] , 
        \input_value[3][124] , \input_value[3][123] , \input_value[3][122] , 
        \input_value[3][121] , \input_value[3][120] , \input_value[3][119] , 
        \input_value[3][118] , \input_value[3][117] , \input_value[3][116] , 
        \input_value[3][115] , \input_value[3][114] , \input_value[3][113] , 
        \input_value[3][112] , \input_value[3][111] , \input_value[3][110] , 
        \input_value[3][109] , \input_value[3][108] , \input_value[3][107] , 
        \input_value[3][106] , \input_value[3][105] , \input_value[3][104] , 
        \input_value[3][103] , \input_value[3][102] , \input_value[3][101] , 
        \input_value[3][100] , \input_value[3][99] , \input_value[3][98] , 
        \input_value[3][97] , \input_value[3][96] , \input_value[3][95] , 
        \input_value[3][94] , \input_value[3][93] , \input_value[3][92] , 
        \input_value[3][91] , \input_value[3][90] , \input_value[3][89] , 
        \input_value[3][88] , \input_value[3][87] , \input_value[3][86] , 
        \input_value[3][85] , \input_value[3][84] , \input_value[3][83] , 
        \input_value[3][82] , \input_value[3][81] , \input_value[3][80] , 
        \input_value[3][79] , \input_value[3][78] , \input_value[3][77] , 
        \input_value[3][76] , \input_value[3][75] , \input_value[3][74] , 
        \input_value[3][73] , \input_value[3][72] , \input_value[3][71] , 
        \input_value[3][70] , \input_value[3][69] , \input_value[3][68] , 
        \input_value[3][67] , \input_value[3][66] , \input_value[3][65] , 
        \input_value[3][64] , \input_value[3][63] , \input_value[3][62] , 
        \input_value[3][61] , \input_value[3][60] , \input_value[3][59] , 
        \input_value[3][58] , \input_value[3][57] , \input_value[3][56] , 
        \input_value[3][55] , \input_value[3][54] , \input_value[3][53] , 
        \input_value[3][52] , \input_value[3][51] , \input_value[3][50] , 
        \input_value[3][49] , \input_value[3][48] , \input_value[3][47] , 
        \input_value[3][46] , \input_value[3][45] , \input_value[3][44] , 
        \input_value[3][43] , \input_value[3][42] , \input_value[3][41] , 
        \input_value[3][40] , \input_value[3][39] , \input_value[3][38] , 
        \input_value[3][37] , \input_value[3][36] , \input_value[3][35] , 
        \input_value[3][34] , \input_value[3][33] , \input_value[3][32] , 
        \input_value[3][31] , \input_value[3][30] , \input_value[3][29] , 
        \input_value[3][28] , \input_value[3][27] , \input_value[3][26] , 
        \input_value[3][25] , \input_value[3][24] , \input_value[3][23] , 
        \input_value[3][22] , \input_value[3][21] , \input_value[3][20] , 
        \input_value[3][19] , \input_value[3][18] , \input_value[3][17] , 
        \input_value[3][16] , \input_value[3][15] , \input_value[3][14] , 
        \input_value[3][13] , \input_value[3][12] , \input_value[3][11] , 
        \input_value[3][10] , \input_value[3][9] , \input_value[3][8] , 
        \input_value[3][7] , \input_value[3][6] , \input_value[3][5] , 
        \input_value[3][4] , \input_value[3][3] , \input_value[3][2] , 
        \input_value[3][1] , \input_value[3][0] }), .input_weight({
        \input_weight[3][127] , \input_weight[3][126] , \input_weight[3][125] , 
        \input_weight[3][124] , \input_weight[3][123] , \input_weight[3][122] , 
        \input_weight[3][121] , \input_weight[3][120] , \input_weight[3][119] , 
        \input_weight[3][118] , \input_weight[3][117] , \input_weight[3][116] , 
        \input_weight[3][115] , \input_weight[3][114] , \input_weight[3][113] , 
        \input_weight[3][112] , \input_weight[3][111] , \input_weight[3][110] , 
        \input_weight[3][109] , \input_weight[3][108] , \input_weight[3][107] , 
        \input_weight[3][106] , \input_weight[3][105] , \input_weight[3][104] , 
        \input_weight[3][103] , \input_weight[3][102] , \input_weight[3][101] , 
        \input_weight[3][100] , \input_weight[3][99] , \input_weight[3][98] , 
        \input_weight[3][97] , \input_weight[3][96] , \input_weight[3][95] , 
        \input_weight[3][94] , \input_weight[3][93] , \input_weight[3][92] , 
        \input_weight[3][91] , \input_weight[3][90] , \input_weight[3][89] , 
        \input_weight[3][88] , \input_weight[3][87] , \input_weight[3][86] , 
        \input_weight[3][85] , \input_weight[3][84] , \input_weight[3][83] , 
        \input_weight[3][82] , \input_weight[3][81] , \input_weight[3][80] , 
        \input_weight[3][79] , \input_weight[3][78] , \input_weight[3][77] , 
        \input_weight[3][76] , \input_weight[3][75] , \input_weight[3][74] , 
        \input_weight[3][73] , \input_weight[3][72] , \input_weight[3][71] , 
        \input_weight[3][70] , \input_weight[3][69] , \input_weight[3][68] , 
        \input_weight[3][67] , \input_weight[3][66] , \input_weight[3][65] , 
        \input_weight[3][64] , \input_weight[3][63] , \input_weight[3][62] , 
        \input_weight[3][61] , \input_weight[3][60] , \input_weight[3][59] , 
        \input_weight[3][58] , \input_weight[3][57] , \input_weight[3][56] , 
        \input_weight[3][55] , \input_weight[3][54] , \input_weight[3][53] , 
        \input_weight[3][52] , \input_weight[3][51] , \input_weight[3][50] , 
        \input_weight[3][49] , \input_weight[3][48] , \input_weight[3][47] , 
        \input_weight[3][46] , \input_weight[3][45] , \input_weight[3][44] , 
        \input_weight[3][43] , \input_weight[3][42] , \input_weight[3][41] , 
        \input_weight[3][40] , \input_weight[3][39] , \input_weight[3][38] , 
        \input_weight[3][37] , \input_weight[3][36] , \input_weight[3][35] , 
        \input_weight[3][34] , \input_weight[3][33] , \input_weight[3][32] , 
        \input_weight[3][31] , \input_weight[3][30] , \input_weight[3][29] , 
        \input_weight[3][28] , \input_weight[3][27] , \input_weight[3][26] , 
        \input_weight[3][25] , \input_weight[3][24] , \input_weight[3][23] , 
        \input_weight[3][22] , \input_weight[3][21] , \input_weight[3][20] , 
        \input_weight[3][19] , \input_weight[3][18] , \input_weight[3][17] , 
        \input_weight[3][16] , \input_weight[3][15] , \input_weight[3][14] , 
        \input_weight[3][13] , \input_weight[3][12] , \input_weight[3][11] , 
        \input_weight[3][10] , \input_weight[3][9] , \input_weight[3][8] , 
        \input_weight[3][7] , \input_weight[3][6] , \input_weight[3][5] , 
        \input_weight[3][4] , \input_weight[3][3] , \input_weight[3][2] , 
        \input_weight[3][1] , \input_weight[3][0] }), .input_bias({
        \input_bias[3][15] , \input_bias[3][14] , \input_bias[3][13] , 
        \input_bias[3][12] , \input_bias[3][11] , \input_bias[3][10] , 
        \input_bias[3][9] , \input_bias[3][8] , \input_bias[3][7] , 
        \input_bias[3][6] , \input_bias[3][5] , \input_bias[3][4] , 
        \input_bias[3][3] , \input_bias[3][2] , \input_bias[3][1] , 
        \input_bias[3][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[3][15] , \output_value[3][14] , \output_value[3][13] , 
        \output_value[3][12] , \output_value[3][11] , \output_value[3][10] , 
        \output_value[3][9] , \output_value[3][8] , \output_value[3][7] , 
        \output_value[3][6] , \output_value[3][5] , \output_value[3][4] , 
        \output_value[3][3] , \output_value[3][2] , \output_value[3][1] , 
        \output_value[3][0] }), .clk(WE) );
  neuron_4 \generate_neurons[4].u_neuron  ( .input_value({
        \input_value[4][127] , \input_value[4][126] , \input_value[4][125] , 
        \input_value[4][124] , \input_value[4][123] , \input_value[4][122] , 
        \input_value[4][121] , \input_value[4][120] , \input_value[4][119] , 
        \input_value[4][118] , \input_value[4][117] , \input_value[4][116] , 
        \input_value[4][115] , \input_value[4][114] , \input_value[4][113] , 
        \input_value[4][112] , \input_value[4][111] , \input_value[4][110] , 
        \input_value[4][109] , \input_value[4][108] , \input_value[4][107] , 
        \input_value[4][106] , \input_value[4][105] , \input_value[4][104] , 
        \input_value[4][103] , \input_value[4][102] , \input_value[4][101] , 
        \input_value[4][100] , \input_value[4][99] , \input_value[4][98] , 
        \input_value[4][97] , \input_value[4][96] , \input_value[4][95] , 
        \input_value[4][94] , \input_value[4][93] , \input_value[4][92] , 
        \input_value[4][91] , \input_value[4][90] , \input_value[4][89] , 
        \input_value[4][88] , \input_value[4][87] , \input_value[4][86] , 
        \input_value[4][85] , \input_value[4][84] , \input_value[4][83] , 
        \input_value[4][82] , \input_value[4][81] , \input_value[4][80] , 
        \input_value[4][79] , \input_value[4][78] , \input_value[4][77] , 
        \input_value[4][76] , \input_value[4][75] , \input_value[4][74] , 
        \input_value[4][73] , \input_value[4][72] , \input_value[4][71] , 
        \input_value[4][70] , \input_value[4][69] , \input_value[4][68] , 
        \input_value[4][67] , \input_value[4][66] , \input_value[4][65] , 
        \input_value[4][64] , \input_value[4][63] , \input_value[4][62] , 
        \input_value[4][61] , \input_value[4][60] , \input_value[4][59] , 
        \input_value[4][58] , \input_value[4][57] , \input_value[4][56] , 
        \input_value[4][55] , \input_value[4][54] , \input_value[4][53] , 
        \input_value[4][52] , \input_value[4][51] , \input_value[4][50] , 
        \input_value[4][49] , \input_value[4][48] , \input_value[4][47] , 
        \input_value[4][46] , \input_value[4][45] , \input_value[4][44] , 
        \input_value[4][43] , \input_value[4][42] , \input_value[4][41] , 
        \input_value[4][40] , \input_value[4][39] , \input_value[4][38] , 
        \input_value[4][37] , \input_value[4][36] , \input_value[4][35] , 
        \input_value[4][34] , \input_value[4][33] , \input_value[4][32] , 
        \input_value[4][31] , \input_value[4][30] , \input_value[4][29] , 
        \input_value[4][28] , \input_value[4][27] , \input_value[4][26] , 
        \input_value[4][25] , \input_value[4][24] , \input_value[4][23] , 
        \input_value[4][22] , \input_value[4][21] , \input_value[4][20] , 
        \input_value[4][19] , \input_value[4][18] , \input_value[4][17] , 
        \input_value[4][16] , \input_value[4][15] , \input_value[4][14] , 
        \input_value[4][13] , \input_value[4][12] , \input_value[4][11] , 
        \input_value[4][10] , \input_value[4][9] , \input_value[4][8] , 
        \input_value[4][7] , \input_value[4][6] , \input_value[4][5] , 
        \input_value[4][4] , \input_value[4][3] , \input_value[4][2] , 
        \input_value[4][1] , \input_value[4][0] }), .input_weight({
        \input_weight[4][127] , \input_weight[4][126] , \input_weight[4][125] , 
        \input_weight[4][124] , \input_weight[4][123] , \input_weight[4][122] , 
        \input_weight[4][121] , \input_weight[4][120] , \input_weight[4][119] , 
        \input_weight[4][118] , \input_weight[4][117] , \input_weight[4][116] , 
        \input_weight[4][115] , \input_weight[4][114] , \input_weight[4][113] , 
        \input_weight[4][112] , \input_weight[4][111] , \input_weight[4][110] , 
        \input_weight[4][109] , \input_weight[4][108] , \input_weight[4][107] , 
        \input_weight[4][106] , \input_weight[4][105] , \input_weight[4][104] , 
        \input_weight[4][103] , \input_weight[4][102] , \input_weight[4][101] , 
        \input_weight[4][100] , \input_weight[4][99] , \input_weight[4][98] , 
        \input_weight[4][97] , \input_weight[4][96] , \input_weight[4][95] , 
        \input_weight[4][94] , \input_weight[4][93] , \input_weight[4][92] , 
        \input_weight[4][91] , \input_weight[4][90] , \input_weight[4][89] , 
        \input_weight[4][88] , \input_weight[4][87] , \input_weight[4][86] , 
        \input_weight[4][85] , \input_weight[4][84] , \input_weight[4][83] , 
        \input_weight[4][82] , \input_weight[4][81] , \input_weight[4][80] , 
        \input_weight[4][79] , \input_weight[4][78] , \input_weight[4][77] , 
        \input_weight[4][76] , \input_weight[4][75] , \input_weight[4][74] , 
        \input_weight[4][73] , \input_weight[4][72] , \input_weight[4][71] , 
        \input_weight[4][70] , \input_weight[4][69] , \input_weight[4][68] , 
        \input_weight[4][67] , \input_weight[4][66] , \input_weight[4][65] , 
        \input_weight[4][64] , \input_weight[4][63] , \input_weight[4][62] , 
        \input_weight[4][61] , \input_weight[4][60] , \input_weight[4][59] , 
        \input_weight[4][58] , \input_weight[4][57] , \input_weight[4][56] , 
        \input_weight[4][55] , \input_weight[4][54] , \input_weight[4][53] , 
        \input_weight[4][52] , \input_weight[4][51] , \input_weight[4][50] , 
        \input_weight[4][49] , \input_weight[4][48] , \input_weight[4][47] , 
        \input_weight[4][46] , \input_weight[4][45] , \input_weight[4][44] , 
        \input_weight[4][43] , \input_weight[4][42] , \input_weight[4][41] , 
        \input_weight[4][40] , \input_weight[4][39] , \input_weight[4][38] , 
        \input_weight[4][37] , \input_weight[4][36] , \input_weight[4][35] , 
        \input_weight[4][34] , \input_weight[4][33] , \input_weight[4][32] , 
        \input_weight[4][31] , \input_weight[4][30] , \input_weight[4][29] , 
        \input_weight[4][28] , \input_weight[4][27] , \input_weight[4][26] , 
        \input_weight[4][25] , \input_weight[4][24] , \input_weight[4][23] , 
        \input_weight[4][22] , \input_weight[4][21] , \input_weight[4][20] , 
        \input_weight[4][19] , \input_weight[4][18] , \input_weight[4][17] , 
        \input_weight[4][16] , \input_weight[4][15] , \input_weight[4][14] , 
        \input_weight[4][13] , \input_weight[4][12] , \input_weight[4][11] , 
        \input_weight[4][10] , \input_weight[4][9] , \input_weight[4][8] , 
        \input_weight[4][7] , \input_weight[4][6] , \input_weight[4][5] , 
        \input_weight[4][4] , \input_weight[4][3] , \input_weight[4][2] , 
        \input_weight[4][1] , \input_weight[4][0] }), .input_bias({
        \input_bias[4][15] , \input_bias[4][14] , \input_bias[4][13] , 
        \input_bias[4][12] , \input_bias[4][11] , \input_bias[4][10] , 
        \input_bias[4][9] , \input_bias[4][8] , \input_bias[4][7] , 
        \input_bias[4][6] , \input_bias[4][5] , \input_bias[4][4] , 
        \input_bias[4][3] , \input_bias[4][2] , \input_bias[4][1] , 
        \input_bias[4][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[4][15] , \output_value[4][14] , \output_value[4][13] , 
        \output_value[4][12] , \output_value[4][11] , \output_value[4][10] , 
        \output_value[4][9] , \output_value[4][8] , \output_value[4][7] , 
        \output_value[4][6] , \output_value[4][5] , \output_value[4][4] , 
        \output_value[4][3] , \output_value[4][2] , \output_value[4][1] , 
        \output_value[4][0] }), .clk(WE) );
  neuron_3 \generate_neurons[5].u_neuron  ( .input_value({
        \input_value[5][127] , \input_value[5][126] , \input_value[5][125] , 
        \input_value[5][124] , \input_value[5][123] , \input_value[5][122] , 
        \input_value[5][121] , \input_value[5][120] , \input_value[5][119] , 
        \input_value[5][118] , \input_value[5][117] , \input_value[5][116] , 
        \input_value[5][115] , \input_value[5][114] , \input_value[5][113] , 
        \input_value[5][112] , \input_value[5][111] , \input_value[5][110] , 
        \input_value[5][109] , \input_value[5][108] , \input_value[5][107] , 
        \input_value[5][106] , \input_value[5][105] , \input_value[5][104] , 
        \input_value[5][103] , \input_value[5][102] , \input_value[5][101] , 
        \input_value[5][100] , \input_value[5][99] , \input_value[5][98] , 
        \input_value[5][97] , \input_value[5][96] , \input_value[5][95] , 
        \input_value[5][94] , \input_value[5][93] , \input_value[5][92] , 
        \input_value[5][91] , \input_value[5][90] , \input_value[5][89] , 
        \input_value[5][88] , \input_value[5][87] , \input_value[5][86] , 
        \input_value[5][85] , \input_value[5][84] , \input_value[5][83] , 
        \input_value[5][82] , \input_value[5][81] , \input_value[5][80] , 
        \input_value[5][79] , \input_value[5][78] , \input_value[5][77] , 
        \input_value[5][76] , \input_value[5][75] , \input_value[5][74] , 
        \input_value[5][73] , \input_value[5][72] , \input_value[5][71] , 
        \input_value[5][70] , \input_value[5][69] , \input_value[5][68] , 
        \input_value[5][67] , \input_value[5][66] , \input_value[5][65] , 
        \input_value[5][64] , \input_value[5][63] , \input_value[5][62] , 
        \input_value[5][61] , \input_value[5][60] , \input_value[5][59] , 
        \input_value[5][58] , \input_value[5][57] , \input_value[5][56] , 
        \input_value[5][55] , \input_value[5][54] , \input_value[5][53] , 
        \input_value[5][52] , \input_value[5][51] , \input_value[5][50] , 
        \input_value[5][49] , \input_value[5][48] , \input_value[5][47] , 
        \input_value[5][46] , \input_value[5][45] , \input_value[5][44] , 
        \input_value[5][43] , \input_value[5][42] , \input_value[5][41] , 
        \input_value[5][40] , \input_value[5][39] , \input_value[5][38] , 
        \input_value[5][37] , \input_value[5][36] , \input_value[5][35] , 
        \input_value[5][34] , \input_value[5][33] , \input_value[5][32] , 
        \input_value[5][31] , \input_value[5][30] , \input_value[5][29] , 
        \input_value[5][28] , \input_value[5][27] , \input_value[5][26] , 
        \input_value[5][25] , \input_value[5][24] , \input_value[5][23] , 
        \input_value[5][22] , \input_value[5][21] , \input_value[5][20] , 
        \input_value[5][19] , \input_value[5][18] , \input_value[5][17] , 
        \input_value[5][16] , \input_value[5][15] , \input_value[5][14] , 
        \input_value[5][13] , \input_value[5][12] , \input_value[5][11] , 
        \input_value[5][10] , \input_value[5][9] , \input_value[5][8] , 
        \input_value[5][7] , \input_value[5][6] , \input_value[5][5] , 
        \input_value[5][4] , \input_value[5][3] , \input_value[5][2] , 
        \input_value[5][1] , \input_value[5][0] }), .input_weight({
        \input_weight[5][127] , \input_weight[5][126] , \input_weight[5][125] , 
        \input_weight[5][124] , \input_weight[5][123] , \input_weight[5][122] , 
        \input_weight[5][121] , \input_weight[5][120] , \input_weight[5][119] , 
        \input_weight[5][118] , \input_weight[5][117] , \input_weight[5][116] , 
        \input_weight[5][115] , \input_weight[5][114] , \input_weight[5][113] , 
        \input_weight[5][112] , \input_weight[5][111] , \input_weight[5][110] , 
        \input_weight[5][109] , \input_weight[5][108] , \input_weight[5][107] , 
        \input_weight[5][106] , \input_weight[5][105] , \input_weight[5][104] , 
        \input_weight[5][103] , \input_weight[5][102] , \input_weight[5][101] , 
        \input_weight[5][100] , \input_weight[5][99] , \input_weight[5][98] , 
        \input_weight[5][97] , \input_weight[5][96] , \input_weight[5][95] , 
        \input_weight[5][94] , \input_weight[5][93] , \input_weight[5][92] , 
        \input_weight[5][91] , \input_weight[5][90] , \input_weight[5][89] , 
        \input_weight[5][88] , \input_weight[5][87] , \input_weight[5][86] , 
        \input_weight[5][85] , \input_weight[5][84] , \input_weight[5][83] , 
        \input_weight[5][82] , \input_weight[5][81] , \input_weight[5][80] , 
        \input_weight[5][79] , \input_weight[5][78] , \input_weight[5][77] , 
        \input_weight[5][76] , \input_weight[5][75] , \input_weight[5][74] , 
        \input_weight[5][73] , \input_weight[5][72] , \input_weight[5][71] , 
        \input_weight[5][70] , \input_weight[5][69] , \input_weight[5][68] , 
        \input_weight[5][67] , \input_weight[5][66] , \input_weight[5][65] , 
        \input_weight[5][64] , \input_weight[5][63] , \input_weight[5][62] , 
        \input_weight[5][61] , \input_weight[5][60] , \input_weight[5][59] , 
        \input_weight[5][58] , \input_weight[5][57] , \input_weight[5][56] , 
        \input_weight[5][55] , \input_weight[5][54] , \input_weight[5][53] , 
        \input_weight[5][52] , \input_weight[5][51] , \input_weight[5][50] , 
        \input_weight[5][49] , \input_weight[5][48] , \input_weight[5][47] , 
        \input_weight[5][46] , \input_weight[5][45] , \input_weight[5][44] , 
        \input_weight[5][43] , \input_weight[5][42] , \input_weight[5][41] , 
        \input_weight[5][40] , \input_weight[5][39] , \input_weight[5][38] , 
        \input_weight[5][37] , \input_weight[5][36] , \input_weight[5][35] , 
        \input_weight[5][34] , \input_weight[5][33] , \input_weight[5][32] , 
        \input_weight[5][31] , \input_weight[5][30] , \input_weight[5][29] , 
        \input_weight[5][28] , \input_weight[5][27] , \input_weight[5][26] , 
        \input_weight[5][25] , \input_weight[5][24] , \input_weight[5][23] , 
        \input_weight[5][22] , \input_weight[5][21] , \input_weight[5][20] , 
        \input_weight[5][19] , \input_weight[5][18] , \input_weight[5][17] , 
        \input_weight[5][16] , \input_weight[5][15] , \input_weight[5][14] , 
        \input_weight[5][13] , \input_weight[5][12] , \input_weight[5][11] , 
        \input_weight[5][10] , \input_weight[5][9] , \input_weight[5][8] , 
        \input_weight[5][7] , \input_weight[5][6] , \input_weight[5][5] , 
        \input_weight[5][4] , \input_weight[5][3] , \input_weight[5][2] , 
        \input_weight[5][1] , \input_weight[5][0] }), .input_bias({
        \input_bias[5][15] , \input_bias[5][14] , \input_bias[5][13] , 
        \input_bias[5][12] , \input_bias[5][11] , \input_bias[5][10] , 
        \input_bias[5][9] , \input_bias[5][8] , \input_bias[5][7] , 
        \input_bias[5][6] , \input_bias[5][5] , \input_bias[5][4] , 
        \input_bias[5][3] , \input_bias[5][2] , \input_bias[5][1] , 
        \input_bias[5][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[5][15] , \output_value[5][14] , \output_value[5][13] , 
        \output_value[5][12] , \output_value[5][11] , \output_value[5][10] , 
        \output_value[5][9] , \output_value[5][8] , \output_value[5][7] , 
        \output_value[5][6] , \output_value[5][5] , \output_value[5][4] , 
        \output_value[5][3] , \output_value[5][2] , \output_value[5][1] , 
        \output_value[5][0] }), .clk(WE) );
  neuron_2 \generate_neurons[6].u_neuron  ( .input_value({
        \input_value[6][127] , \input_value[6][126] , \input_value[6][125] , 
        \input_value[6][124] , \input_value[6][123] , \input_value[6][122] , 
        \input_value[6][121] , \input_value[6][120] , \input_value[6][119] , 
        \input_value[6][118] , \input_value[6][117] , \input_value[6][116] , 
        \input_value[6][115] , \input_value[6][114] , \input_value[6][113] , 
        \input_value[6][112] , \input_value[6][111] , \input_value[6][110] , 
        \input_value[6][109] , \input_value[6][108] , \input_value[6][107] , 
        \input_value[6][106] , \input_value[6][105] , \input_value[6][104] , 
        \input_value[6][103] , \input_value[6][102] , \input_value[6][101] , 
        \input_value[6][100] , \input_value[6][99] , \input_value[6][98] , 
        \input_value[6][97] , \input_value[6][96] , \input_value[6][95] , 
        \input_value[6][94] , \input_value[6][93] , \input_value[6][92] , 
        \input_value[6][91] , \input_value[6][90] , \input_value[6][89] , 
        \input_value[6][88] , \input_value[6][87] , \input_value[6][86] , 
        \input_value[6][85] , \input_value[6][84] , \input_value[6][83] , 
        \input_value[6][82] , \input_value[6][81] , \input_value[6][80] , 
        \input_value[6][79] , \input_value[6][78] , \input_value[6][77] , 
        \input_value[6][76] , \input_value[6][75] , \input_value[6][74] , 
        \input_value[6][73] , \input_value[6][72] , \input_value[6][71] , 
        \input_value[6][70] , \input_value[6][69] , \input_value[6][68] , 
        \input_value[6][67] , \input_value[6][66] , \input_value[6][65] , 
        \input_value[6][64] , \input_value[6][63] , \input_value[6][62] , 
        \input_value[6][61] , \input_value[6][60] , \input_value[6][59] , 
        \input_value[6][58] , \input_value[6][57] , \input_value[6][56] , 
        \input_value[6][55] , \input_value[6][54] , \input_value[6][53] , 
        \input_value[6][52] , \input_value[6][51] , \input_value[6][50] , 
        \input_value[6][49] , \input_value[6][48] , \input_value[6][47] , 
        \input_value[6][46] , \input_value[6][45] , \input_value[6][44] , 
        \input_value[6][43] , \input_value[6][42] , \input_value[6][41] , 
        \input_value[6][40] , \input_value[6][39] , \input_value[6][38] , 
        \input_value[6][37] , \input_value[6][36] , \input_value[6][35] , 
        \input_value[6][34] , \input_value[6][33] , \input_value[6][32] , 
        \input_value[6][31] , \input_value[6][30] , \input_value[6][29] , 
        \input_value[6][28] , \input_value[6][27] , \input_value[6][26] , 
        \input_value[6][25] , \input_value[6][24] , \input_value[6][23] , 
        \input_value[6][22] , \input_value[6][21] , \input_value[6][20] , 
        \input_value[6][19] , \input_value[6][18] , \input_value[6][17] , 
        \input_value[6][16] , \input_value[6][15] , \input_value[6][14] , 
        \input_value[6][13] , \input_value[6][12] , \input_value[6][11] , 
        \input_value[6][10] , \input_value[6][9] , \input_value[6][8] , 
        \input_value[6][7] , \input_value[6][6] , \input_value[6][5] , 
        \input_value[6][4] , \input_value[6][3] , \input_value[6][2] , 
        \input_value[6][1] , \input_value[6][0] }), .input_weight({
        \input_weight[6][127] , \input_weight[6][126] , \input_weight[6][125] , 
        \input_weight[6][124] , \input_weight[6][123] , \input_weight[6][122] , 
        \input_weight[6][121] , \input_weight[6][120] , \input_weight[6][119] , 
        \input_weight[6][118] , \input_weight[6][117] , \input_weight[6][116] , 
        \input_weight[6][115] , \input_weight[6][114] , \input_weight[6][113] , 
        \input_weight[6][112] , \input_weight[6][111] , \input_weight[6][110] , 
        \input_weight[6][109] , \input_weight[6][108] , \input_weight[6][107] , 
        \input_weight[6][106] , \input_weight[6][105] , \input_weight[6][104] , 
        \input_weight[6][103] , \input_weight[6][102] , \input_weight[6][101] , 
        \input_weight[6][100] , \input_weight[6][99] , \input_weight[6][98] , 
        \input_weight[6][97] , \input_weight[6][96] , \input_weight[6][95] , 
        \input_weight[6][94] , \input_weight[6][93] , \input_weight[6][92] , 
        \input_weight[6][91] , \input_weight[6][90] , \input_weight[6][89] , 
        \input_weight[6][88] , \input_weight[6][87] , \input_weight[6][86] , 
        \input_weight[6][85] , \input_weight[6][84] , \input_weight[6][83] , 
        \input_weight[6][82] , \input_weight[6][81] , \input_weight[6][80] , 
        \input_weight[6][79] , \input_weight[6][78] , \input_weight[6][77] , 
        \input_weight[6][76] , \input_weight[6][75] , \input_weight[6][74] , 
        \input_weight[6][73] , \input_weight[6][72] , \input_weight[6][71] , 
        \input_weight[6][70] , \input_weight[6][69] , \input_weight[6][68] , 
        \input_weight[6][67] , \input_weight[6][66] , \input_weight[6][65] , 
        \input_weight[6][64] , \input_weight[6][63] , \input_weight[6][62] , 
        \input_weight[6][61] , \input_weight[6][60] , \input_weight[6][59] , 
        \input_weight[6][58] , \input_weight[6][57] , \input_weight[6][56] , 
        \input_weight[6][55] , \input_weight[6][54] , \input_weight[6][53] , 
        \input_weight[6][52] , \input_weight[6][51] , \input_weight[6][50] , 
        \input_weight[6][49] , \input_weight[6][48] , \input_weight[6][47] , 
        \input_weight[6][46] , \input_weight[6][45] , \input_weight[6][44] , 
        \input_weight[6][43] , \input_weight[6][42] , \input_weight[6][41] , 
        \input_weight[6][40] , \input_weight[6][39] , \input_weight[6][38] , 
        \input_weight[6][37] , \input_weight[6][36] , \input_weight[6][35] , 
        \input_weight[6][34] , \input_weight[6][33] , \input_weight[6][32] , 
        \input_weight[6][31] , \input_weight[6][30] , \input_weight[6][29] , 
        \input_weight[6][28] , \input_weight[6][27] , \input_weight[6][26] , 
        \input_weight[6][25] , \input_weight[6][24] , \input_weight[6][23] , 
        \input_weight[6][22] , \input_weight[6][21] , \input_weight[6][20] , 
        \input_weight[6][19] , \input_weight[6][18] , \input_weight[6][17] , 
        \input_weight[6][16] , \input_weight[6][15] , \input_weight[6][14] , 
        \input_weight[6][13] , \input_weight[6][12] , \input_weight[6][11] , 
        \input_weight[6][10] , \input_weight[6][9] , \input_weight[6][8] , 
        \input_weight[6][7] , \input_weight[6][6] , \input_weight[6][5] , 
        \input_weight[6][4] , \input_weight[6][3] , \input_weight[6][2] , 
        \input_weight[6][1] , \input_weight[6][0] }), .input_bias({
        \input_bias[6][15] , \input_bias[6][14] , \input_bias[6][13] , 
        \input_bias[6][12] , \input_bias[6][11] , \input_bias[6][10] , 
        \input_bias[6][9] , \input_bias[6][8] , \input_bias[6][7] , 
        \input_bias[6][6] , \input_bias[6][5] , \input_bias[6][4] , 
        \input_bias[6][3] , \input_bias[6][2] , \input_bias[6][1] , 
        \input_bias[6][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[6][15] , \output_value[6][14] , \output_value[6][13] , 
        \output_value[6][12] , \output_value[6][11] , \output_value[6][10] , 
        \output_value[6][9] , \output_value[6][8] , \output_value[6][7] , 
        \output_value[6][6] , \output_value[6][5] , \output_value[6][4] , 
        \output_value[6][3] , \output_value[6][2] , \output_value[6][1] , 
        \output_value[6][0] }), .clk(WE) );
  neuron_1 \generate_neurons[7].u_neuron  ( .input_value({
        \input_value[7][127] , \input_value[7][126] , \input_value[7][125] , 
        \input_value[7][124] , \input_value[7][123] , \input_value[7][122] , 
        \input_value[7][121] , \input_value[7][120] , \input_value[7][119] , 
        \input_value[7][118] , \input_value[7][117] , \input_value[7][116] , 
        \input_value[7][115] , \input_value[7][114] , \input_value[7][113] , 
        \input_value[7][112] , \input_value[7][111] , \input_value[7][110] , 
        \input_value[7][109] , \input_value[7][108] , \input_value[7][107] , 
        \input_value[7][106] , \input_value[7][105] , \input_value[7][104] , 
        \input_value[7][103] , \input_value[7][102] , \input_value[7][101] , 
        \input_value[7][100] , \input_value[7][99] , \input_value[7][98] , 
        \input_value[7][97] , \input_value[7][96] , \input_value[7][95] , 
        \input_value[7][94] , \input_value[7][93] , \input_value[7][92] , 
        \input_value[7][91] , \input_value[7][90] , \input_value[7][89] , 
        \input_value[7][88] , \input_value[7][87] , \input_value[7][86] , 
        \input_value[7][85] , \input_value[7][84] , \input_value[7][83] , 
        \input_value[7][82] , \input_value[7][81] , \input_value[7][80] , 
        \input_value[7][79] , \input_value[7][78] , \input_value[7][77] , 
        \input_value[7][76] , \input_value[7][75] , \input_value[7][74] , 
        \input_value[7][73] , \input_value[7][72] , \input_value[7][71] , 
        \input_value[7][70] , \input_value[7][69] , \input_value[7][68] , 
        \input_value[7][67] , \input_value[7][66] , \input_value[7][65] , 
        \input_value[7][64] , \input_value[7][63] , \input_value[7][62] , 
        \input_value[7][61] , \input_value[7][60] , \input_value[7][59] , 
        \input_value[7][58] , \input_value[7][57] , \input_value[7][56] , 
        \input_value[7][55] , \input_value[7][54] , \input_value[7][53] , 
        \input_value[7][52] , \input_value[7][51] , \input_value[7][50] , 
        \input_value[7][49] , \input_value[7][48] , \input_value[7][47] , 
        \input_value[7][46] , \input_value[7][45] , \input_value[7][44] , 
        \input_value[7][43] , \input_value[7][42] , \input_value[7][41] , 
        \input_value[7][40] , \input_value[7][39] , \input_value[7][38] , 
        \input_value[7][37] , \input_value[7][36] , \input_value[7][35] , 
        \input_value[7][34] , \input_value[7][33] , \input_value[7][32] , 
        \input_value[7][31] , \input_value[7][30] , \input_value[7][29] , 
        \input_value[7][28] , \input_value[7][27] , \input_value[7][26] , 
        \input_value[7][25] , \input_value[7][24] , \input_value[7][23] , 
        \input_value[7][22] , \input_value[7][21] , \input_value[7][20] , 
        \input_value[7][19] , \input_value[7][18] , \input_value[7][17] , 
        \input_value[7][16] , \input_value[7][15] , \input_value[7][14] , 
        \input_value[7][13] , \input_value[7][12] , \input_value[7][11] , 
        \input_value[7][10] , \input_value[7][9] , \input_value[7][8] , 
        \input_value[7][7] , \input_value[7][6] , \input_value[7][5] , 
        \input_value[7][4] , \input_value[7][3] , \input_value[7][2] , 
        \input_value[7][1] , \input_value[7][0] }), .input_weight({
        \input_weight[7][127] , \input_weight[7][126] , \input_weight[7][125] , 
        \input_weight[7][124] , \input_weight[7][123] , \input_weight[7][122] , 
        \input_weight[7][121] , \input_weight[7][120] , \input_weight[7][119] , 
        \input_weight[7][118] , \input_weight[7][117] , \input_weight[7][116] , 
        \input_weight[7][115] , \input_weight[7][114] , \input_weight[7][113] , 
        \input_weight[7][112] , \input_weight[7][111] , \input_weight[7][110] , 
        \input_weight[7][109] , \input_weight[7][108] , \input_weight[7][107] , 
        \input_weight[7][106] , \input_weight[7][105] , \input_weight[7][104] , 
        \input_weight[7][103] , \input_weight[7][102] , \input_weight[7][101] , 
        \input_weight[7][100] , \input_weight[7][99] , \input_weight[7][98] , 
        \input_weight[7][97] , \input_weight[7][96] , \input_weight[7][95] , 
        \input_weight[7][94] , \input_weight[7][93] , \input_weight[7][92] , 
        \input_weight[7][91] , \input_weight[7][90] , \input_weight[7][89] , 
        \input_weight[7][88] , \input_weight[7][87] , \input_weight[7][86] , 
        \input_weight[7][85] , \input_weight[7][84] , \input_weight[7][83] , 
        \input_weight[7][82] , \input_weight[7][81] , \input_weight[7][80] , 
        \input_weight[7][79] , \input_weight[7][78] , \input_weight[7][77] , 
        \input_weight[7][76] , \input_weight[7][75] , \input_weight[7][74] , 
        \input_weight[7][73] , \input_weight[7][72] , \input_weight[7][71] , 
        \input_weight[7][70] , \input_weight[7][69] , \input_weight[7][68] , 
        \input_weight[7][67] , \input_weight[7][66] , \input_weight[7][65] , 
        \input_weight[7][64] , \input_weight[7][63] , \input_weight[7][62] , 
        \input_weight[7][61] , \input_weight[7][60] , \input_weight[7][59] , 
        \input_weight[7][58] , \input_weight[7][57] , \input_weight[7][56] , 
        \input_weight[7][55] , \input_weight[7][54] , \input_weight[7][53] , 
        \input_weight[7][52] , \input_weight[7][51] , \input_weight[7][50] , 
        \input_weight[7][49] , \input_weight[7][48] , \input_weight[7][47] , 
        \input_weight[7][46] , \input_weight[7][45] , \input_weight[7][44] , 
        \input_weight[7][43] , \input_weight[7][42] , \input_weight[7][41] , 
        \input_weight[7][40] , \input_weight[7][39] , \input_weight[7][38] , 
        \input_weight[7][37] , \input_weight[7][36] , \input_weight[7][35] , 
        \input_weight[7][34] , \input_weight[7][33] , \input_weight[7][32] , 
        \input_weight[7][31] , \input_weight[7][30] , \input_weight[7][29] , 
        \input_weight[7][28] , \input_weight[7][27] , \input_weight[7][26] , 
        \input_weight[7][25] , \input_weight[7][24] , \input_weight[7][23] , 
        \input_weight[7][22] , \input_weight[7][21] , \input_weight[7][20] , 
        \input_weight[7][19] , \input_weight[7][18] , \input_weight[7][17] , 
        \input_weight[7][16] , \input_weight[7][15] , \input_weight[7][14] , 
        \input_weight[7][13] , \input_weight[7][12] , \input_weight[7][11] , 
        \input_weight[7][10] , \input_weight[7][9] , \input_weight[7][8] , 
        \input_weight[7][7] , \input_weight[7][6] , \input_weight[7][5] , 
        \input_weight[7][4] , \input_weight[7][3] , \input_weight[7][2] , 
        \input_weight[7][1] , \input_weight[7][0] }), .input_bias({
        \input_bias[7][15] , \input_bias[7][14] , \input_bias[7][13] , 
        \input_bias[7][12] , \input_bias[7][11] , \input_bias[7][10] , 
        \input_bias[7][9] , \input_bias[7][8] , \input_bias[7][7] , 
        \input_bias[7][6] , \input_bias[7][5] , \input_bias[7][4] , 
        \input_bias[7][3] , \input_bias[7][2] , \input_bias[7][1] , 
        \input_bias[7][0] }), .rst(rst), .en(RE), .srdy(RE), .output_value({
        \output_value[7][15] , \output_value[7][14] , \output_value[7][13] , 
        \output_value[7][12] , \output_value[7][11] , \output_value[7][10] , 
        \output_value[7][9] , \output_value[7][8] , \output_value[7][7] , 
        \output_value[7][6] , \output_value[7][5] , \output_value[7][4] , 
        \output_value[7][3] , \output_value[7][2] , \output_value[7][1] , 
        \output_value[7][0] }), .clk(WE) );
  arbiter u_fwd_arbiter ( .neuron_done({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .rst(rst), .network({\forward_network[7][31] , 
        \forward_network[7][30] , \forward_network[7][29] , 
        \forward_network[7][28] , \forward_network[7][27] , 
        \forward_network[7][26] , \forward_network[7][25] , 
        \forward_network[7][24] , \forward_network[7][23] , 
        \forward_network[7][22] , \forward_network[7][21] , 
        \forward_network[7][20] , \forward_network[7][19] , 
        \forward_network[7][18] , \forward_network[7][17] , 
        \forward_network[7][16] , \forward_network[7][15] , 
        \forward_network[7][14] , \forward_network[7][13] , 
        \forward_network[7][12] , \forward_network[7][11] , 
        \forward_network[7][10] , \forward_network[7][9] , 
        \forward_network[7][8] , \forward_network[7][7] , 
        \forward_network[7][6] , \forward_network[7][5] , 
        \forward_network[7][4] , \forward_network[7][3] , 
        \forward_network[7][2] , \forward_network[7][1] , 
        \forward_network[7][0] , \forward_network[6][31] , 
        \forward_network[6][30] , \forward_network[6][29] , 
        \forward_network[6][28] , \forward_network[6][27] , 
        \forward_network[6][26] , \forward_network[6][25] , 
        \forward_network[6][24] , \forward_network[6][23] , 
        \forward_network[6][22] , \forward_network[6][21] , 
        \forward_network[6][20] , \forward_network[6][19] , 
        \forward_network[6][18] , \forward_network[6][17] , 
        \forward_network[6][16] , \forward_network[6][15] , 
        \forward_network[6][14] , \forward_network[6][13] , 
        \forward_network[6][12] , \forward_network[6][11] , 
        \forward_network[6][10] , \forward_network[6][9] , 
        \forward_network[6][8] , \forward_network[6][7] , 
        \forward_network[6][6] , \forward_network[6][5] , 
        \forward_network[6][4] , \forward_network[6][3] , 
        \forward_network[6][2] , \forward_network[6][1] , 
        \forward_network[6][0] , \forward_network[5][31] , 
        \forward_network[5][30] , \forward_network[5][29] , 
        \forward_network[5][28] , \forward_network[5][27] , 
        \forward_network[5][26] , \forward_network[5][25] , 
        \forward_network[5][24] , \forward_network[5][23] , 
        \forward_network[5][22] , \forward_network[5][21] , 
        \forward_network[5][20] , \forward_network[5][19] , 
        \forward_network[5][18] , \forward_network[5][17] , 
        \forward_network[5][16] , \forward_network[5][15] , 
        \forward_network[5][14] , \forward_network[5][13] , 
        \forward_network[5][12] , \forward_network[5][11] , 
        \forward_network[5][10] , \forward_network[5][9] , 
        \forward_network[5][8] , \forward_network[5][7] , 
        \forward_network[5][6] , \forward_network[5][5] , 
        \forward_network[5][4] , \forward_network[5][3] , 
        \forward_network[5][2] , \forward_network[5][1] , 
        \forward_network[5][0] , \forward_network[4][31] , 
        \forward_network[4][30] , \forward_network[4][29] , 
        \forward_network[4][28] , \forward_network[4][27] , 
        \forward_network[4][26] , \forward_network[4][25] , 
        \forward_network[4][24] , \forward_network[4][23] , 
        \forward_network[4][22] , \forward_network[4][21] , 
        \forward_network[4][20] , \forward_network[4][19] , 
        \forward_network[4][18] , \forward_network[4][17] , 
        \forward_network[4][16] , \forward_network[4][15] , 
        \forward_network[4][14] , \forward_network[4][13] , 
        \forward_network[4][12] , \forward_network[4][11] , 
        \forward_network[4][10] , \forward_network[4][9] , 
        \forward_network[4][8] , \forward_network[4][7] , 
        \forward_network[4][6] , \forward_network[4][5] , 
        \forward_network[4][4] , \forward_network[4][3] , 
        \forward_network[4][2] , \forward_network[4][1] , 
        \forward_network[4][0] , \forward_network[3][31] , 
        \forward_network[3][30] , \forward_network[3][29] , 
        \forward_network[3][28] , \forward_network[3][27] , 
        \forward_network[3][26] , \forward_network[3][25] , 
        \forward_network[3][24] , \forward_network[3][23] , 
        \forward_network[3][22] , \forward_network[3][21] , 
        \forward_network[3][20] , \forward_network[3][19] , 
        \forward_network[3][18] , \forward_network[3][17] , 
        \forward_network[3][16] , \forward_network[3][15] , 
        \forward_network[3][14] , \forward_network[3][13] , 
        \forward_network[3][12] , \forward_network[3][11] , 
        \forward_network[3][10] , \forward_network[3][9] , 
        \forward_network[3][8] , \forward_network[3][7] , 
        \forward_network[3][6] , \forward_network[3][5] , 
        \forward_network[3][4] , \forward_network[3][3] , 
        \forward_network[3][2] , \forward_network[3][1] , 
        \forward_network[3][0] , \forward_network[2][31] , 
        \forward_network[2][30] , \forward_network[2][29] , 
        \forward_network[2][28] , \forward_network[2][27] , 
        \forward_network[2][26] , \forward_network[2][25] , 
        \forward_network[2][24] , \forward_network[2][23] , 
        \forward_network[2][22] , \forward_network[2][21] , 
        \forward_network[2][20] , \forward_network[2][19] , 
        \forward_network[2][18] , \forward_network[2][17] , 
        \forward_network[2][16] , \forward_network[2][15] , 
        \forward_network[2][14] , \forward_network[2][13] , 
        \forward_network[2][12] , \forward_network[2][11] , 
        \forward_network[2][10] , \forward_network[2][9] , 
        \forward_network[2][8] , \forward_network[2][7] , 
        \forward_network[2][6] , \forward_network[2][5] , 
        \forward_network[2][4] , \forward_network[2][3] , 
        \forward_network[2][2] , \forward_network[2][1] , 
        \forward_network[2][0] , \forward_network[1][31] , 
        \forward_network[1][30] , \forward_network[1][29] , 
        \forward_network[1][28] , \forward_network[1][27] , 
        \forward_network[1][26] , \forward_network[1][25] , 
        \forward_network[1][24] , \forward_network[1][23] , 
        \forward_network[1][22] , \forward_network[1][21] , 
        \forward_network[1][20] , \forward_network[1][19] , 
        \forward_network[1][18] , \forward_network[1][17] , 
        \forward_network[1][16] , \forward_network[1][15] , 
        \forward_network[1][14] , \forward_network[1][13] , 
        \forward_network[1][12] , \forward_network[1][11] , 
        \forward_network[1][10] , \forward_network[1][9] , 
        \forward_network[1][8] , \forward_network[1][7] , 
        \forward_network[1][6] , \forward_network[1][5] , 
        \forward_network[1][4] , \forward_network[1][3] , 
        \forward_network[1][2] , \forward_network[1][1] , 
        \forward_network[1][0] , \forward_network[0][31] , 
        \forward_network[0][30] , \forward_network[0][29] , 
        \forward_network[0][28] , \forward_network[0][27] , 
        \forward_network[0][26] , \forward_network[0][25] , 
        \forward_network[0][24] , \forward_network[0][23] , 
        \forward_network[0][22] , \forward_network[0][21] , 
        \forward_network[0][20] , \forward_network[0][19] , 
        \forward_network[0][18] , \forward_network[0][17] , 
        \forward_network[0][16] , \forward_network[0][15] , 
        \forward_network[0][14] , \forward_network[0][13] , 
        \forward_network[0][12] , \forward_network[0][11] , 
        \forward_network[0][10] , \forward_network[0][9] , 
        \forward_network[0][8] , \forward_network[0][7] , 
        \forward_network[0][6] , \forward_network[0][5] , 
        \forward_network[0][4] , \forward_network[0][3] , 
        \forward_network[0][2] , \forward_network[0][1] , 
        \forward_network[0][0] }) );
  routing_engine u_fwd_routing_engine ( .port_dest({WE, WE, WE, WE, WE, WE, WE, 
        WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, WE, 
        WE, WE, WE, WE, WE, WE, WE}), .control({SYNOPSYS_UNCONNECTED__0, 
        fwd_routing_engine_control[18:16], SYNOPSYS_UNCONNECTED__1, 
        fwd_routing_engine_control[14], SYNOPSYS_UNCONNECTED__2, 
        fwd_routing_engine_control[12:0]}) );
  benes u_fwd_benes ( .out_output(layer_data_out), .in_input({
        \output_value[0][15] , \output_value[0][14] , \output_value[0][13] , 
        \output_value[0][12] , \output_value[0][11] , \output_value[0][10] , 
        \output_value[0][9] , \output_value[0][8] , \output_value[0][7] , 
        \output_value[0][6] , \output_value[0][5] , \output_value[0][4] , 
        \output_value[0][3] , \output_value[0][2] , \output_value[0][1] , 
        \output_value[0][0] , \output_value[1][15] , \output_value[1][14] , 
        \output_value[1][13] , \output_value[1][12] , \output_value[1][11] , 
        \output_value[1][10] , \output_value[1][9] , \output_value[1][8] , 
        \output_value[1][7] , \output_value[1][6] , \output_value[1][5] , 
        \output_value[1][4] , \output_value[1][3] , \output_value[1][2] , 
        \output_value[1][1] , \output_value[1][0] , \output_value[2][15] , 
        \output_value[2][14] , \output_value[2][13] , \output_value[2][12] , 
        \output_value[2][11] , \output_value[2][10] , \output_value[2][9] , 
        \output_value[2][8] , \output_value[2][7] , \output_value[2][6] , 
        \output_value[2][5] , \output_value[2][4] , \output_value[2][3] , 
        \output_value[2][2] , \output_value[2][1] , \output_value[2][0] , 
        \output_value[3][15] , \output_value[3][14] , \output_value[3][13] , 
        \output_value[3][12] , \output_value[3][11] , \output_value[3][10] , 
        \output_value[3][9] , \output_value[3][8] , \output_value[3][7] , 
        \output_value[3][6] , \output_value[3][5] , \output_value[3][4] , 
        \output_value[3][3] , \output_value[3][2] , \output_value[3][1] , 
        \output_value[3][0] , \output_value[4][15] , \output_value[4][14] , 
        \output_value[4][13] , \output_value[4][12] , \output_value[4][11] , 
        \output_value[4][10] , \output_value[4][9] , \output_value[4][8] , 
        \output_value[4][7] , \output_value[4][6] , \output_value[4][5] , 
        \output_value[4][4] , \output_value[4][3] , \output_value[4][2] , 
        \output_value[4][1] , \output_value[4][0] , \output_value[5][15] , 
        \output_value[5][14] , \output_value[5][13] , \output_value[5][12] , 
        \output_value[5][11] , \output_value[5][10] , \output_value[5][9] , 
        \output_value[5][8] , \output_value[5][7] , \output_value[5][6] , 
        \output_value[5][5] , \output_value[5][4] , \output_value[5][3] , 
        \output_value[5][2] , \output_value[5][1] , \output_value[5][0] , 
        \output_value[6][15] , \output_value[6][14] , \output_value[6][13] , 
        \output_value[6][12] , \output_value[6][11] , \output_value[6][10] , 
        \output_value[6][9] , \output_value[6][8] , \output_value[6][7] , 
        \output_value[6][6] , \output_value[6][5] , \output_value[6][4] , 
        \output_value[6][3] , \output_value[6][2] , \output_value[6][1] , 
        \output_value[6][0] , \output_value[7][15] , \output_value[7][14] , 
        \output_value[7][13] , \output_value[7][12] , \output_value[7][11] , 
        \output_value[7][10] , \output_value[7][9] , \output_value[7][8] , 
        \output_value[7][7] , \output_value[7][6] , \output_value[7][5] , 
        \output_value[7][4] , \output_value[7][3] , \output_value[7][2] , 
        \output_value[7][1] , \output_value[7][0] }), .in_control({1'b0, 
        fwd_routing_engine_control[18:16], 1'b0, 
        fwd_routing_engine_control[14], 1'b0, fwd_routing_engine_control[12:0]}), .port_en_n(1'b1) );
  EDFQD1 \cur_state_reg[2]  ( .D(nxt_state[2]), .E(N156), .CP(clk), .Q(
        cur_state[2]) );
  EDFQD1 \neuron_BAR_reg[5]  ( .D(N115), .E(N114), .CP(clk), .Q(neuron_BAR[5])
         );
  EDFQD1 \neuron_BAR_reg[3]  ( .D(N116), .E(N114), .CP(clk), .Q(neuron_BAR[3])
         );
  EDFQD1 \neuron_BAR_reg[8]  ( .D(N120), .E(N114), .CP(clk), .Q(neuron_BAR[8])
         );
  EDFQD1 \neuron_BAR_reg[6]  ( .D(N118), .E(N114), .CP(clk), .Q(neuron_BAR[6])
         );
  EDFQD1 \neuron_BAR_reg[4]  ( .D(N117), .E(N114), .CP(clk), .Q(neuron_BAR[4])
         );
  EDFQD1 \cur_state_reg[3]  ( .D(nxt_state[3]), .E(N156), .CP(clk), .Q(
        cur_state[3]) );
  EDFQD1 \neuron_BAR_reg[2]  ( .D(N115), .E(N114), .CP(clk), .Q(neuron_BAR[2])
         );
  EDFQD1 \neuron_BAR_reg[7]  ( .D(N119), .E(N114), .CP(clk), .Q(neuron_BAR[7])
         );
  EDFQD1 \neuron_BAR_reg[9]  ( .D(N121), .E(N114), .CP(clk), .Q(neuron_BAR[9])
         );
  EDFQD1 \mem_cur_state_reg[3]  ( .D(mem_nxt_state[3]), .E(N428), .CP(clk), 
        .Q(mem_cur_state[3]) );
  EDFQD1 \mem_cur_state_reg[2]  ( .D(mem_nxt_state[2]), .E(N428), .CP(clk), 
        .Q(mem_cur_state[2]) );
  EDFQD1 \cur_state_reg[1]  ( .D(nxt_state[1]), .E(N156), .CP(clk), .Q(
        cur_state[1]) );
  EDFQD1 \mem_cur_state_reg[1]  ( .D(mem_nxt_state[1]), .E(N428), .CP(clk), 
        .Q(mem_cur_state[1]) );
  EDFQD1 \mem_cur_state_reg[0]  ( .D(mem_nxt_state[0]), .E(N428), .CP(clk), 
        .Q(mem_cur_state[0]) );
  EDFQD1 \cur_state_reg[0]  ( .D(nxt_state[0]), .E(N156), .CP(clk), .Q(
        cur_state[0]) );
  EDFQD1 \nxt_state_reg[0]  ( .D(N123), .E(N122), .CP(clk), .Q(nxt_state[0])
         );
  EDFQD1 \nxt_state_reg[2]  ( .D(N125), .E(N122), .CP(clk), .Q(nxt_state[2])
         );
  EDFQD1 \nxt_state_reg[1]  ( .D(N124), .E(N122), .CP(clk), .Q(nxt_state[1])
         );
  EDFQD1 \nxt_state_reg[3]  ( .D(n585), .E(N122), .CP(clk), .Q(nxt_state[3])
         );
  EDFQD1 \forward_network_reg[4][9]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][9] ) );
  EDFQD1 \forward_network_reg[4][10]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][10] ) );
  EDFQD1 \forward_network_reg[4][11]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][11] ) );
  EDFQD1 \forward_network_reg[4][12]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][12] ) );
  EDFQD1 \forward_network_reg[4][13]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][13] ) );
  EDFQD1 \forward_network_reg[4][14]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][14] ) );
  EDFQD1 \forward_network_reg[4][15]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][15] ) );
  EDFQD1 \forward_network_reg[4][16]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][16] ) );
  EDFQD1 \forward_network_reg[4][17]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][17] ) );
  EDFQD1 \forward_network_reg[4][18]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][18] ) );
  EDFQD1 \forward_network_reg[4][19]  ( .D(WE), .E(n287), .CP(clk), .Q(
        \forward_network[4][19] ) );
  EDFQD1 \forward_network_reg[4][20]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][20] ) );
  EDFQD1 \forward_network_reg[4][21]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][21] ) );
  EDFQD1 \forward_network_reg[4][22]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][22] ) );
  EDFQD1 \forward_network_reg[4][23]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][23] ) );
  EDFQD1 \forward_network_reg[4][24]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][24] ) );
  EDFQD1 \forward_network_reg[4][25]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][25] ) );
  EDFQD1 \forward_network_reg[4][26]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][26] ) );
  EDFQD1 \forward_network_reg[4][27]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][27] ) );
  EDFQD1 \forward_network_reg[4][28]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][28] ) );
  EDFQD1 \forward_network_reg[4][29]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][29] ) );
  EDFQD1 \forward_network_reg[4][30]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][30] ) );
  EDFQD1 \forward_network_reg[4][31]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[4][31] ) );
  EDFQD1 \forward_network_reg[5][9]  ( .D(WE), .E(n286), .CP(clk), .Q(
        \forward_network[5][9] ) );
  EDFQD1 \forward_network_reg[5][10]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][10] ) );
  EDFQD1 \forward_network_reg[5][11]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][11] ) );
  EDFQD1 \forward_network_reg[5][12]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][12] ) );
  EDFQD1 \forward_network_reg[5][13]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][13] ) );
  EDFQD1 \forward_network_reg[5][14]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][14] ) );
  EDFQD1 \forward_network_reg[5][15]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][15] ) );
  EDFQD1 \forward_network_reg[5][16]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][16] ) );
  EDFQD1 \forward_network_reg[5][17]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][17] ) );
  EDFQD1 \forward_network_reg[5][18]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][18] ) );
  EDFQD1 \forward_network_reg[5][19]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][19] ) );
  EDFQD1 \forward_network_reg[5][20]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][20] ) );
  EDFQD1 \forward_network_reg[5][21]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][21] ) );
  EDFQD1 \forward_network_reg[5][22]  ( .D(WE), .E(n285), .CP(clk), .Q(
        \forward_network[5][22] ) );
  EDFQD1 \forward_network_reg[5][23]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][23] ) );
  EDFQD1 \forward_network_reg[5][24]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][24] ) );
  EDFQD1 \forward_network_reg[5][25]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][25] ) );
  EDFQD1 \forward_network_reg[5][26]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][26] ) );
  EDFQD1 \forward_network_reg[5][27]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][27] ) );
  EDFQD1 \forward_network_reg[5][28]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][28] ) );
  EDFQD1 \forward_network_reg[5][29]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][29] ) );
  EDFQD1 \forward_network_reg[5][30]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][30] ) );
  EDFQD1 \forward_network_reg[5][31]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[5][31] ) );
  EDFQD1 \forward_network_reg[6][9]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[6][9] ) );
  EDFQD1 \forward_network_reg[6][10]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[6][10] ) );
  EDFQD1 \forward_network_reg[6][11]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[6][11] ) );
  EDFQD1 \forward_network_reg[6][12]  ( .D(WE), .E(n284), .CP(clk), .Q(
        \forward_network[6][12] ) );
  EDFQD1 \forward_network_reg[6][13]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][13] ) );
  EDFQD1 \forward_network_reg[6][14]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][14] ) );
  EDFQD1 \forward_network_reg[6][15]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][15] ) );
  EDFQD1 \forward_network_reg[6][16]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][16] ) );
  EDFQD1 \forward_network_reg[6][17]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][17] ) );
  EDFQD1 \forward_network_reg[6][18]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][18] ) );
  EDFQD1 \forward_network_reg[6][19]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][19] ) );
  EDFQD1 \forward_network_reg[6][20]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][20] ) );
  EDFQD1 \forward_network_reg[6][21]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][21] ) );
  EDFQD1 \forward_network_reg[6][22]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][22] ) );
  EDFQD1 \forward_network_reg[6][23]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][23] ) );
  EDFQD1 \forward_network_reg[6][24]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][24] ) );
  EDFQD1 \forward_network_reg[6][25]  ( .D(WE), .E(n283), .CP(clk), .Q(
        \forward_network[6][25] ) );
  EDFQD1 \forward_network_reg[6][26]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][26] ) );
  EDFQD1 \forward_network_reg[6][27]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][27] ) );
  EDFQD1 \forward_network_reg[6][28]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][28] ) );
  EDFQD1 \forward_network_reg[6][29]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][29] ) );
  EDFQD1 \forward_network_reg[6][30]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][30] ) );
  EDFQD1 \forward_network_reg[6][31]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[6][31] ) );
  EDFQD1 \forward_network_reg[7][31]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][31] ) );
  EDFQD1 \forward_network_reg[7][30]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][30] ) );
  EDFQD1 \forward_network_reg[7][29]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][29] ) );
  EDFQD1 \forward_network_reg[7][28]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][28] ) );
  EDFQD1 \forward_network_reg[7][27]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][27] ) );
  EDFQD1 \forward_network_reg[7][26]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][26] ) );
  EDFQD1 \forward_network_reg[7][25]  ( .D(WE), .E(n282), .CP(clk), .Q(
        \forward_network[7][25] ) );
  EDFQD1 \forward_network_reg[7][24]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][24] ) );
  EDFQD1 \forward_network_reg[7][23]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][23] ) );
  EDFQD1 \forward_network_reg[7][22]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][22] ) );
  EDFQD1 \forward_network_reg[7][21]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][21] ) );
  EDFQD1 \forward_network_reg[7][20]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][20] ) );
  EDFQD1 \forward_network_reg[7][19]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][19] ) );
  EDFQD1 \forward_network_reg[7][18]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][18] ) );
  EDFQD1 \forward_network_reg[7][17]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][17] ) );
  EDFQD1 \forward_network_reg[7][16]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][16] ) );
  EDFQD1 \forward_network_reg[7][15]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][15] ) );
  EDFQD1 \forward_network_reg[7][14]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][14] ) );
  EDFQD1 \forward_network_reg[7][13]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][13] ) );
  EDFQD1 \forward_network_reg[7][12]  ( .D(WE), .E(n281), .CP(clk), .Q(
        \forward_network[7][12] ) );
  EDFQD1 \forward_network_reg[7][11]  ( .D(WE), .E(n280), .CP(clk), .Q(
        \forward_network[7][11] ) );
  EDFQD1 \forward_network_reg[7][10]  ( .D(WE), .E(n280), .CP(clk), .Q(
        \forward_network[7][10] ) );
  EDFQD1 \forward_network_reg[7][9]  ( .D(WE), .E(n280), .CP(clk), .Q(
        \forward_network[7][9] ) );
  EDFQD1 \forward_network_reg[0][9]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][9] ) );
  EDFQD1 \forward_network_reg[0][10]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][10] ) );
  EDFQD1 \forward_network_reg[0][11]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][11] ) );
  EDFQD1 \forward_network_reg[0][12]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][12] ) );
  EDFQD1 \forward_network_reg[0][13]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][13] ) );
  EDFQD1 \forward_network_reg[0][14]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][14] ) );
  EDFQD1 \forward_network_reg[0][15]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][15] ) );
  EDFQD1 \forward_network_reg[0][16]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][16] ) );
  EDFQD1 \forward_network_reg[0][17]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][17] ) );
  EDFQD1 \forward_network_reg[0][18]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][18] ) );
  EDFQD1 \forward_network_reg[0][19]  ( .D(WE), .E(n272), .CP(clk), .Q(
        \forward_network[0][19] ) );
  EDFQD1 \forward_network_reg[0][20]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][20] ) );
  EDFQD1 \forward_network_reg[0][21]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][21] ) );
  EDFQD1 \forward_network_reg[0][22]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][22] ) );
  EDFQD1 \forward_network_reg[0][23]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][23] ) );
  EDFQD1 \forward_network_reg[0][24]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][24] ) );
  EDFQD1 \forward_network_reg[0][25]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][25] ) );
  EDFQD1 \forward_network_reg[0][26]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][26] ) );
  EDFQD1 \forward_network_reg[0][27]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][27] ) );
  EDFQD1 \forward_network_reg[0][28]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][28] ) );
  EDFQD1 \forward_network_reg[0][29]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][29] ) );
  EDFQD1 \forward_network_reg[0][30]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][30] ) );
  EDFQD1 \forward_network_reg[0][31]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[0][31] ) );
  EDFQD1 \forward_network_reg[1][9]  ( .D(WE), .E(n271), .CP(clk), .Q(
        \forward_network[1][9] ) );
  EDFQD1 \forward_network_reg[1][10]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][10] ) );
  EDFQD1 \forward_network_reg[1][11]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][11] ) );
  EDFQD1 \forward_network_reg[1][12]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][12] ) );
  EDFQD1 \forward_network_reg[1][13]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][13] ) );
  EDFQD1 \forward_network_reg[1][14]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][14] ) );
  EDFQD1 \forward_network_reg[1][15]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][15] ) );
  EDFQD1 \forward_network_reg[1][16]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][16] ) );
  EDFQD1 \forward_network_reg[1][17]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][17] ) );
  EDFQD1 \forward_network_reg[1][18]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][18] ) );
  EDFQD1 \forward_network_reg[1][19]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][19] ) );
  EDFQD1 \forward_network_reg[1][20]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][20] ) );
  EDFQD1 \forward_network_reg[1][21]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][21] ) );
  EDFQD1 \forward_network_reg[1][22]  ( .D(WE), .E(n270), .CP(clk), .Q(
        \forward_network[1][22] ) );
  EDFQD1 \forward_network_reg[1][23]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][23] ) );
  EDFQD1 \forward_network_reg[1][24]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][24] ) );
  EDFQD1 \forward_network_reg[1][25]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][25] ) );
  EDFQD1 \forward_network_reg[1][26]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][26] ) );
  EDFQD1 \forward_network_reg[1][27]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][27] ) );
  EDFQD1 \forward_network_reg[1][28]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][28] ) );
  EDFQD1 \forward_network_reg[1][29]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][29] ) );
  EDFQD1 \forward_network_reg[1][30]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][30] ) );
  EDFQD1 \forward_network_reg[1][31]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[1][31] ) );
  EDFQD1 \forward_network_reg[2][9]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[2][9] ) );
  EDFQD1 \forward_network_reg[2][10]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[2][10] ) );
  EDFQD1 \forward_network_reg[2][11]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[2][11] ) );
  EDFQD1 \forward_network_reg[2][12]  ( .D(WE), .E(n269), .CP(clk), .Q(
        \forward_network[2][12] ) );
  EDFQD1 \forward_network_reg[2][13]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][13] ) );
  EDFQD1 \forward_network_reg[2][14]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][14] ) );
  EDFQD1 \forward_network_reg[2][15]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][15] ) );
  EDFQD1 \forward_network_reg[2][16]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][16] ) );
  EDFQD1 \forward_network_reg[2][17]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][17] ) );
  EDFQD1 \forward_network_reg[2][18]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][18] ) );
  EDFQD1 \forward_network_reg[2][19]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][19] ) );
  EDFQD1 \forward_network_reg[2][20]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][20] ) );
  EDFQD1 \forward_network_reg[2][21]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][21] ) );
  EDFQD1 \forward_network_reg[2][22]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][22] ) );
  EDFQD1 \forward_network_reg[2][23]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][23] ) );
  EDFQD1 \forward_network_reg[2][24]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][24] ) );
  EDFQD1 \forward_network_reg[2][25]  ( .D(WE), .E(n268), .CP(clk), .Q(
        \forward_network[2][25] ) );
  EDFQD1 \forward_network_reg[2][26]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][26] ) );
  EDFQD1 \forward_network_reg[2][27]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][27] ) );
  EDFQD1 \forward_network_reg[2][28]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][28] ) );
  EDFQD1 \forward_network_reg[2][29]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][29] ) );
  EDFQD1 \forward_network_reg[2][30]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][30] ) );
  EDFQD1 \forward_network_reg[2][31]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[2][31] ) );
  EDFQD1 \forward_network_reg[3][31]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][31] ) );
  EDFQD1 \forward_network_reg[3][30]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][30] ) );
  EDFQD1 \forward_network_reg[3][29]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][29] ) );
  EDFQD1 \forward_network_reg[3][28]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][28] ) );
  EDFQD1 \forward_network_reg[3][27]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][27] ) );
  EDFQD1 \forward_network_reg[3][26]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][26] ) );
  EDFQD1 \forward_network_reg[3][25]  ( .D(WE), .E(n267), .CP(clk), .Q(
        \forward_network[3][25] ) );
  EDFQD1 \forward_network_reg[3][24]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][24] ) );
  EDFQD1 \forward_network_reg[3][23]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][23] ) );
  EDFQD1 \forward_network_reg[3][22]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][22] ) );
  EDFQD1 \forward_network_reg[3][21]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][21] ) );
  EDFQD1 \forward_network_reg[3][20]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][20] ) );
  EDFQD1 \forward_network_reg[3][19]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][19] ) );
  EDFQD1 \forward_network_reg[3][18]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][18] ) );
  EDFQD1 \forward_network_reg[3][17]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][17] ) );
  EDFQD1 \forward_network_reg[3][16]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][16] ) );
  EDFQD1 \forward_network_reg[3][15]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][15] ) );
  EDFQD1 \forward_network_reg[3][14]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][14] ) );
  EDFQD1 \forward_network_reg[3][13]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][13] ) );
  EDFQD1 \forward_network_reg[3][12]  ( .D(WE), .E(n266), .CP(clk), .Q(
        \forward_network[3][12] ) );
  EDFQD1 \forward_network_reg[3][11]  ( .D(WE), .E(n265), .CP(clk), .Q(
        \forward_network[3][11] ) );
  EDFQD1 \forward_network_reg[3][10]  ( .D(WE), .E(n265), .CP(clk), .Q(
        \forward_network[3][10] ) );
  EDFQD1 \forward_network_reg[3][9]  ( .D(WE), .E(n265), .CP(clk), .Q(
        \forward_network[3][9] ) );
  EDFQD1 \forward_network_reg[4][0]  ( .D(data_in[95]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][0] ) );
  EDFQD1 \forward_network_reg[4][1]  ( .D(data_in[96]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][1] ) );
  EDFQD1 \forward_network_reg[4][2]  ( .D(data_in[97]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][2] ) );
  EDFQD1 \forward_network_reg[4][3]  ( .D(data_in[98]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][3] ) );
  EDFQD1 \forward_network_reg[4][4]  ( .D(data_in[99]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][4] ) );
  EDFQD1 \forward_network_reg[4][5]  ( .D(data_in[100]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][5] ) );
  EDFQD1 \forward_network_reg[4][6]  ( .D(data_in[101]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][6] ) );
  EDFQD1 \forward_network_reg[4][7]  ( .D(data_in[102]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][7] ) );
  EDFQD1 \forward_network_reg[4][8]  ( .D(data_in[103]), .E(n278), .CP(clk), 
        .Q(\forward_network[4][8] ) );
  EDFQD1 \forward_network_reg[5][0]  ( .D(data_in[103]), .E(n278), .CP(clk), 
        .Q(\forward_network[5][0] ) );
  EDFQD1 \forward_network_reg[5][1]  ( .D(data_in[104]), .E(n278), .CP(clk), 
        .Q(\forward_network[5][1] ) );
  EDFQD1 \forward_network_reg[5][2]  ( .D(data_in[105]), .E(n278), .CP(clk), 
        .Q(\forward_network[5][2] ) );
  EDFQD1 \forward_network_reg[5][3]  ( .D(data_in[106]), .E(n278), .CP(clk), 
        .Q(\forward_network[5][3] ) );
  EDFQD1 \forward_network_reg[5][4]  ( .D(data_in[107]), .E(n279), .CP(clk), 
        .Q(\forward_network[5][4] ) );
  EDFQD1 \forward_network_reg[5][5]  ( .D(data_in[108]), .E(n279), .CP(clk), 
        .Q(\forward_network[5][5] ) );
  EDFQD1 \forward_network_reg[5][6]  ( .D(data_in[109]), .E(n279), .CP(clk), 
        .Q(\forward_network[5][6] ) );
  EDFQD1 \forward_network_reg[5][7]  ( .D(data_in[110]), .E(n279), .CP(clk), 
        .Q(\forward_network[5][7] ) );
  EDFQD1 \forward_network_reg[5][8]  ( .D(data_in[111]), .E(n279), .CP(clk), 
        .Q(\forward_network[5][8] ) );
  EDFQD1 \forward_network_reg[6][0]  ( .D(data_in[111]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][0] ) );
  EDFQD1 \forward_network_reg[6][1]  ( .D(data_in[112]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][1] ) );
  EDFQD1 \forward_network_reg[6][2]  ( .D(data_in[113]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][2] ) );
  EDFQD1 \forward_network_reg[6][3]  ( .D(data_in[114]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][3] ) );
  EDFQD1 \forward_network_reg[6][4]  ( .D(data_in[115]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][4] ) );
  EDFQD1 \forward_network_reg[6][5]  ( .D(data_in[116]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][5] ) );
  EDFQD1 \forward_network_reg[6][6]  ( .D(data_in[117]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][6] ) );
  EDFQD1 \forward_network_reg[6][7]  ( .D(data_in[118]), .E(n279), .CP(clk), 
        .Q(\forward_network[6][7] ) );
  EDFQD1 \forward_network_reg[6][8]  ( .D(data_in[119]), .E(n280), .CP(clk), 
        .Q(\forward_network[6][8] ) );
  EDFQD1 \forward_network_reg[7][0]  ( .D(data_in[119]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][0] ) );
  EDFQD1 \forward_network_reg[7][1]  ( .D(data_in[120]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][1] ) );
  EDFQD1 \forward_network_reg[7][2]  ( .D(data_in[121]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][2] ) );
  EDFQD1 \forward_network_reg[7][8]  ( .D(data_in[127]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][8] ) );
  EDFQD1 \forward_network_reg[7][7]  ( .D(data_in[126]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][7] ) );
  EDFQD1 \forward_network_reg[7][6]  ( .D(data_in[125]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][6] ) );
  EDFQD1 \forward_network_reg[7][5]  ( .D(data_in[124]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][5] ) );
  EDFQD1 \forward_network_reg[7][4]  ( .D(data_in[123]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][4] ) );
  EDFQD1 \forward_network_reg[7][3]  ( .D(data_in[122]), .E(n280), .CP(clk), 
        .Q(\forward_network[7][3] ) );
  EDFQD1 \forward_network_reg[0][0]  ( .D(data_in[95]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][0] ) );
  EDFQD1 \forward_network_reg[0][1]  ( .D(data_in[96]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][1] ) );
  EDFQD1 \forward_network_reg[0][2]  ( .D(data_in[97]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][2] ) );
  EDFQD1 \forward_network_reg[0][3]  ( .D(data_in[98]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][3] ) );
  EDFQD1 \forward_network_reg[0][4]  ( .D(data_in[99]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][4] ) );
  EDFQD1 \forward_network_reg[0][5]  ( .D(data_in[100]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][5] ) );
  EDFQD1 \forward_network_reg[0][6]  ( .D(data_in[101]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][6] ) );
  EDFQD1 \forward_network_reg[0][7]  ( .D(data_in[102]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][7] ) );
  EDFQD1 \forward_network_reg[0][8]  ( .D(data_in[103]), .E(n263), .CP(clk), 
        .Q(\forward_network[0][8] ) );
  EDFQD1 \forward_network_reg[1][0]  ( .D(data_in[103]), .E(n263), .CP(clk), 
        .Q(\forward_network[1][0] ) );
  EDFQD1 \forward_network_reg[1][1]  ( .D(data_in[104]), .E(n263), .CP(clk), 
        .Q(\forward_network[1][1] ) );
  EDFQD1 \forward_network_reg[1][2]  ( .D(data_in[105]), .E(n263), .CP(clk), 
        .Q(\forward_network[1][2] ) );
  EDFQD1 \forward_network_reg[1][3]  ( .D(data_in[106]), .E(n263), .CP(clk), 
        .Q(\forward_network[1][3] ) );
  EDFQD1 \forward_network_reg[1][4]  ( .D(data_in[107]), .E(n264), .CP(clk), 
        .Q(\forward_network[1][4] ) );
  EDFQD1 \forward_network_reg[1][5]  ( .D(data_in[108]), .E(n264), .CP(clk), 
        .Q(\forward_network[1][5] ) );
  EDFQD1 \forward_network_reg[1][6]  ( .D(data_in[109]), .E(n264), .CP(clk), 
        .Q(\forward_network[1][6] ) );
  EDFQD1 \forward_network_reg[1][7]  ( .D(data_in[110]), .E(n264), .CP(clk), 
        .Q(\forward_network[1][7] ) );
  EDFQD1 \forward_network_reg[1][8]  ( .D(data_in[111]), .E(n264), .CP(clk), 
        .Q(\forward_network[1][8] ) );
  EDFQD1 \forward_network_reg[2][0]  ( .D(data_in[111]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][0] ) );
  EDFQD1 \forward_network_reg[2][1]  ( .D(data_in[112]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][1] ) );
  EDFQD1 \forward_network_reg[2][2]  ( .D(data_in[113]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][2] ) );
  EDFQD1 \forward_network_reg[2][3]  ( .D(data_in[114]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][3] ) );
  EDFQD1 \forward_network_reg[2][4]  ( .D(data_in[115]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][4] ) );
  EDFQD1 \forward_network_reg[2][5]  ( .D(data_in[116]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][5] ) );
  EDFQD1 \forward_network_reg[2][6]  ( .D(data_in[117]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][6] ) );
  EDFQD1 \forward_network_reg[2][7]  ( .D(data_in[118]), .E(n264), .CP(clk), 
        .Q(\forward_network[2][7] ) );
  EDFQD1 \forward_network_reg[2][8]  ( .D(data_in[119]), .E(n265), .CP(clk), 
        .Q(\forward_network[2][8] ) );
  EDFQD1 \forward_network_reg[3][0]  ( .D(data_in[119]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][0] ) );
  EDFQD1 \forward_network_reg[3][1]  ( .D(data_in[120]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][1] ) );
  EDFQD1 \forward_network_reg[3][2]  ( .D(data_in[121]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][2] ) );
  EDFQD1 \forward_network_reg[3][8]  ( .D(data_in[127]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][8] ) );
  EDFQD1 \forward_network_reg[3][7]  ( .D(data_in[126]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][7] ) );
  EDFQD1 \forward_network_reg[3][6]  ( .D(data_in[125]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][6] ) );
  EDFQD1 \forward_network_reg[3][5]  ( .D(data_in[124]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][5] ) );
  EDFQD1 \forward_network_reg[3][4]  ( .D(data_in[123]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][4] ) );
  EDFQD1 \forward_network_reg[3][3]  ( .D(data_in[122]), .E(n265), .CP(clk), 
        .Q(\forward_network[3][3] ) );
  EDFQD1 \input_weight_reg[6][99]  ( .D(data_in[99]), .E(n437), .CP(clk), .Q(
        \input_weight[6][99] ) );
  EDFQD1 \input_weight_reg[6][100]  ( .D(data_in[100]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][100] ) );
  EDFQD1 \input_weight_reg[6][101]  ( .D(data_in[101]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][101] ) );
  EDFQD1 \input_weight_reg[6][102]  ( .D(data_in[102]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][102] ) );
  EDFQD1 \input_weight_reg[6][103]  ( .D(data_in[103]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][103] ) );
  EDFQD1 \input_weight_reg[6][104]  ( .D(data_in[104]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][104] ) );
  EDFQD1 \input_weight_reg[6][105]  ( .D(data_in[105]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][105] ) );
  EDFQD1 \input_weight_reg[6][106]  ( .D(data_in[106]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][106] ) );
  EDFQD1 \input_weight_reg[6][107]  ( .D(data_in[107]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][107] ) );
  EDFQD1 \input_weight_reg[6][108]  ( .D(data_in[108]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][108] ) );
  EDFQD1 \input_weight_reg[6][109]  ( .D(data_in[109]), .E(n437), .CP(clk), 
        .Q(\input_weight[6][109] ) );
  EDFQD1 \input_weight_reg[6][110]  ( .D(data_in[110]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][110] ) );
  EDFQD1 \input_weight_reg[6][111]  ( .D(data_in[111]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][111] ) );
  EDFQD1 \input_weight_reg[6][112]  ( .D(data_in[112]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][112] ) );
  EDFQD1 \input_weight_reg[6][113]  ( .D(data_in[113]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][113] ) );
  EDFQD1 \input_weight_reg[6][114]  ( .D(data_in[114]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][114] ) );
  EDFQD1 \input_weight_reg[6][115]  ( .D(data_in[115]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][115] ) );
  EDFQD1 \input_weight_reg[6][116]  ( .D(data_in[116]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][116] ) );
  EDFQD1 \input_weight_reg[6][117]  ( .D(data_in[117]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][117] ) );
  EDFQD1 \input_weight_reg[6][118]  ( .D(data_in[118]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][118] ) );
  EDFQD1 \input_weight_reg[6][119]  ( .D(data_in[119]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][119] ) );
  EDFQD1 \input_weight_reg[6][120]  ( .D(data_in[120]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][120] ) );
  EDFQD1 \input_weight_reg[6][121]  ( .D(data_in[121]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][121] ) );
  EDFQD1 \input_weight_reg[6][122]  ( .D(data_in[122]), .E(n436), .CP(clk), 
        .Q(\input_weight[6][122] ) );
  EDFQD1 \input_weight_reg[6][123]  ( .D(data_in[123]), .E(n435), .CP(clk), 
        .Q(\input_weight[6][123] ) );
  EDFQD1 \input_weight_reg[6][124]  ( .D(data_in[124]), .E(n435), .CP(clk), 
        .Q(\input_weight[6][124] ) );
  EDFQD1 \input_weight_reg[6][125]  ( .D(data_in[125]), .E(n435), .CP(clk), 
        .Q(\input_weight[6][125] ) );
  EDFQD1 \input_weight_reg[6][126]  ( .D(data_in[126]), .E(n435), .CP(clk), 
        .Q(\input_weight[6][126] ) );
  EDFQD1 \input_weight_reg[6][127]  ( .D(data_in[127]), .E(n435), .CP(clk), 
        .Q(\input_weight[6][127] ) );
  EDFQD1 \input_weight_reg[6][98]  ( .D(data_in[98]), .E(n435), .CP(clk), .Q(
        \input_weight[6][98] ) );
  EDFQD1 \input_weight_reg[6][97]  ( .D(data_in[97]), .E(n435), .CP(clk), .Q(
        \input_weight[6][97] ) );
  EDFQD1 \input_weight_reg[6][96]  ( .D(data_in[96]), .E(n435), .CP(clk), .Q(
        \input_weight[6][96] ) );
  EDFQD1 \input_weight_reg[6][95]  ( .D(data_in[95]), .E(n435), .CP(clk), .Q(
        \input_weight[6][95] ) );
  EDFQD1 \input_weight_reg[6][94]  ( .D(data_in[94]), .E(n435), .CP(clk), .Q(
        \input_weight[6][94] ) );
  EDFQD1 \input_weight_reg[6][93]  ( .D(data_in[93]), .E(n435), .CP(clk), .Q(
        \input_weight[6][93] ) );
  EDFQD1 \input_weight_reg[6][92]  ( .D(data_in[92]), .E(n435), .CP(clk), .Q(
        \input_weight[6][92] ) );
  EDFQD1 \input_weight_reg[6][91]  ( .D(data_in[91]), .E(n435), .CP(clk), .Q(
        \input_weight[6][91] ) );
  EDFQD1 \input_weight_reg[6][90]  ( .D(data_in[90]), .E(n434), .CP(clk), .Q(
        \input_weight[6][90] ) );
  EDFQD1 \input_weight_reg[6][89]  ( .D(data_in[89]), .E(n434), .CP(clk), .Q(
        \input_weight[6][89] ) );
  EDFQD1 \input_weight_reg[6][88]  ( .D(data_in[88]), .E(n434), .CP(clk), .Q(
        \input_weight[6][88] ) );
  EDFQD1 \input_weight_reg[6][87]  ( .D(data_in[87]), .E(n434), .CP(clk), .Q(
        \input_weight[6][87] ) );
  EDFQD1 \input_weight_reg[6][86]  ( .D(data_in[86]), .E(n434), .CP(clk), .Q(
        \input_weight[6][86] ) );
  EDFQD1 \input_weight_reg[6][85]  ( .D(data_in[85]), .E(n434), .CP(clk), .Q(
        \input_weight[6][85] ) );
  EDFQD1 \input_weight_reg[6][84]  ( .D(data_in[84]), .E(n434), .CP(clk), .Q(
        \input_weight[6][84] ) );
  EDFQD1 \input_weight_reg[6][83]  ( .D(data_in[83]), .E(n434), .CP(clk), .Q(
        \input_weight[6][83] ) );
  EDFQD1 \input_weight_reg[6][82]  ( .D(data_in[82]), .E(n434), .CP(clk), .Q(
        \input_weight[6][82] ) );
  EDFQD1 \input_weight_reg[6][81]  ( .D(data_in[81]), .E(n434), .CP(clk), .Q(
        \input_weight[6][81] ) );
  EDFQD1 \input_weight_reg[6][80]  ( .D(data_in[80]), .E(n434), .CP(clk), .Q(
        \input_weight[6][80] ) );
  EDFQD1 \input_weight_reg[6][79]  ( .D(data_in[79]), .E(n434), .CP(clk), .Q(
        \input_weight[6][79] ) );
  EDFQD1 \input_weight_reg[6][78]  ( .D(data_in[78]), .E(n434), .CP(clk), .Q(
        \input_weight[6][78] ) );
  EDFQD1 \input_weight_reg[6][77]  ( .D(data_in[77]), .E(n433), .CP(clk), .Q(
        \input_weight[6][77] ) );
  EDFQD1 \input_weight_reg[6][76]  ( .D(data_in[76]), .E(n433), .CP(clk), .Q(
        \input_weight[6][76] ) );
  EDFQD1 \input_weight_reg[6][75]  ( .D(data_in[75]), .E(n433), .CP(clk), .Q(
        \input_weight[6][75] ) );
  EDFQD1 \input_weight_reg[6][74]  ( .D(data_in[74]), .E(n433), .CP(clk), .Q(
        \input_weight[6][74] ) );
  EDFQD1 \input_weight_reg[6][73]  ( .D(data_in[73]), .E(n433), .CP(clk), .Q(
        \input_weight[6][73] ) );
  EDFQD1 \input_weight_reg[6][72]  ( .D(data_in[72]), .E(n433), .CP(clk), .Q(
        \input_weight[6][72] ) );
  EDFQD1 \input_weight_reg[6][71]  ( .D(data_in[71]), .E(n433), .CP(clk), .Q(
        \input_weight[6][71] ) );
  EDFQD1 \input_weight_reg[6][70]  ( .D(data_in[70]), .E(n433), .CP(clk), .Q(
        \input_weight[6][70] ) );
  EDFQD1 \input_weight_reg[6][69]  ( .D(data_in[69]), .E(n433), .CP(clk), .Q(
        \input_weight[6][69] ) );
  EDFQD1 \input_weight_reg[6][68]  ( .D(data_in[68]), .E(n433), .CP(clk), .Q(
        \input_weight[6][68] ) );
  EDFQD1 \input_weight_reg[6][67]  ( .D(data_in[67]), .E(n433), .CP(clk), .Q(
        \input_weight[6][67] ) );
  EDFQD1 \input_weight_reg[6][66]  ( .D(data_in[66]), .E(n433), .CP(clk), .Q(
        \input_weight[6][66] ) );
  EDFQD1 \input_weight_reg[6][65]  ( .D(data_in[65]), .E(n433), .CP(clk), .Q(
        \input_weight[6][65] ) );
  EDFQD1 \input_weight_reg[6][64]  ( .D(data_in[64]), .E(n432), .CP(clk), .Q(
        \input_weight[6][64] ) );
  EDFQD1 \input_weight_reg[6][63]  ( .D(data_in[63]), .E(n432), .CP(clk), .Q(
        \input_weight[6][63] ) );
  EDFQD1 \input_weight_reg[6][62]  ( .D(data_in[62]), .E(n432), .CP(clk), .Q(
        \input_weight[6][62] ) );
  EDFQD1 \input_weight_reg[6][61]  ( .D(data_in[61]), .E(n432), .CP(clk), .Q(
        \input_weight[6][61] ) );
  EDFQD1 \input_weight_reg[6][60]  ( .D(data_in[60]), .E(n432), .CP(clk), .Q(
        \input_weight[6][60] ) );
  EDFQD1 \input_weight_reg[6][59]  ( .D(data_in[59]), .E(n432), .CP(clk), .Q(
        \input_weight[6][59] ) );
  EDFQD1 \input_weight_reg[6][58]  ( .D(data_in[58]), .E(n432), .CP(clk), .Q(
        \input_weight[6][58] ) );
  EDFQD1 \input_weight_reg[6][57]  ( .D(data_in[57]), .E(n432), .CP(clk), .Q(
        \input_weight[6][57] ) );
  EDFQD1 \input_weight_reg[6][56]  ( .D(data_in[56]), .E(n432), .CP(clk), .Q(
        \input_weight[6][56] ) );
  EDFQD1 \input_weight_reg[6][55]  ( .D(data_in[55]), .E(n432), .CP(clk), .Q(
        \input_weight[6][55] ) );
  EDFQD1 \input_weight_reg[6][54]  ( .D(data_in[54]), .E(n432), .CP(clk), .Q(
        \input_weight[6][54] ) );
  EDFQD1 \input_weight_reg[6][53]  ( .D(data_in[53]), .E(n432), .CP(clk), .Q(
        \input_weight[6][53] ) );
  EDFQD1 \input_weight_reg[6][52]  ( .D(data_in[52]), .E(n432), .CP(clk), .Q(
        \input_weight[6][52] ) );
  EDFQD1 \input_weight_reg[6][51]  ( .D(data_in[51]), .E(n431), .CP(clk), .Q(
        \input_weight[6][51] ) );
  EDFQD1 \input_weight_reg[6][50]  ( .D(data_in[50]), .E(n431), .CP(clk), .Q(
        \input_weight[6][50] ) );
  EDFQD1 \input_weight_reg[6][49]  ( .D(data_in[49]), .E(n431), .CP(clk), .Q(
        \input_weight[6][49] ) );
  EDFQD1 \input_weight_reg[6][48]  ( .D(data_in[48]), .E(n431), .CP(clk), .Q(
        \input_weight[6][48] ) );
  EDFQD1 \input_weight_reg[6][47]  ( .D(data_in[47]), .E(n431), .CP(clk), .Q(
        \input_weight[6][47] ) );
  EDFQD1 \input_weight_reg[6][46]  ( .D(data_in[46]), .E(n431), .CP(clk), .Q(
        \input_weight[6][46] ) );
  EDFQD1 \input_weight_reg[6][45]  ( .D(data_in[45]), .E(n431), .CP(clk), .Q(
        \input_weight[6][45] ) );
  EDFQD1 \input_weight_reg[6][44]  ( .D(data_in[44]), .E(n431), .CP(clk), .Q(
        \input_weight[6][44] ) );
  EDFQD1 \input_weight_reg[6][43]  ( .D(data_in[43]), .E(n431), .CP(clk), .Q(
        \input_weight[6][43] ) );
  EDFQD1 \input_weight_reg[6][42]  ( .D(data_in[42]), .E(n431), .CP(clk), .Q(
        \input_weight[6][42] ) );
  EDFQD1 \input_weight_reg[6][41]  ( .D(data_in[41]), .E(n431), .CP(clk), .Q(
        \input_weight[6][41] ) );
  EDFQD1 \input_weight_reg[6][40]  ( .D(data_in[40]), .E(n431), .CP(clk), .Q(
        \input_weight[6][40] ) );
  EDFQD1 \input_weight_reg[6][39]  ( .D(data_in[39]), .E(n431), .CP(clk), .Q(
        \input_weight[6][39] ) );
  EDFQD1 \input_weight_reg[6][38]  ( .D(data_in[38]), .E(n430), .CP(clk), .Q(
        \input_weight[6][38] ) );
  EDFQD1 \input_weight_reg[6][37]  ( .D(data_in[37]), .E(n430), .CP(clk), .Q(
        \input_weight[6][37] ) );
  EDFQD1 \input_weight_reg[6][36]  ( .D(data_in[36]), .E(n430), .CP(clk), .Q(
        \input_weight[6][36] ) );
  EDFQD1 \input_weight_reg[6][35]  ( .D(data_in[35]), .E(n430), .CP(clk), .Q(
        \input_weight[6][35] ) );
  EDFQD1 \input_weight_reg[6][34]  ( .D(data_in[34]), .E(n430), .CP(clk), .Q(
        \input_weight[6][34] ) );
  EDFQD1 \input_weight_reg[6][33]  ( .D(data_in[33]), .E(n430), .CP(clk), .Q(
        \input_weight[6][33] ) );
  EDFQD1 \input_weight_reg[6][32]  ( .D(data_in[32]), .E(n430), .CP(clk), .Q(
        \input_weight[6][32] ) );
  EDFQD1 \input_weight_reg[6][31]  ( .D(data_in[31]), .E(n430), .CP(clk), .Q(
        \input_weight[6][31] ) );
  EDFQD1 \input_weight_reg[6][30]  ( .D(data_in[30]), .E(n430), .CP(clk), .Q(
        \input_weight[6][30] ) );
  EDFQD1 \input_weight_reg[6][29]  ( .D(data_in[29]), .E(n430), .CP(clk), .Q(
        \input_weight[6][29] ) );
  EDFQD1 \input_weight_reg[6][28]  ( .D(data_in[28]), .E(n430), .CP(clk), .Q(
        \input_weight[6][28] ) );
  EDFQD1 \input_weight_reg[6][27]  ( .D(data_in[27]), .E(n430), .CP(clk), .Q(
        \input_weight[6][27] ) );
  EDFQD1 \input_weight_reg[6][26]  ( .D(data_in[26]), .E(n430), .CP(clk), .Q(
        \input_weight[6][26] ) );
  EDFQD1 \input_weight_reg[6][25]  ( .D(data_in[25]), .E(n429), .CP(clk), .Q(
        \input_weight[6][25] ) );
  EDFQD1 \input_weight_reg[6][24]  ( .D(data_in[24]), .E(n429), .CP(clk), .Q(
        \input_weight[6][24] ) );
  EDFQD1 \input_weight_reg[6][23]  ( .D(data_in[23]), .E(n429), .CP(clk), .Q(
        \input_weight[6][23] ) );
  EDFQD1 \input_weight_reg[6][22]  ( .D(data_in[22]), .E(n429), .CP(clk), .Q(
        \input_weight[6][22] ) );
  EDFQD1 \input_weight_reg[6][21]  ( .D(data_in[21]), .E(n429), .CP(clk), .Q(
        \input_weight[6][21] ) );
  EDFQD1 \input_weight_reg[6][20]  ( .D(data_in[20]), .E(n429), .CP(clk), .Q(
        \input_weight[6][20] ) );
  EDFQD1 \input_weight_reg[6][19]  ( .D(data_in[19]), .E(n429), .CP(clk), .Q(
        \input_weight[6][19] ) );
  EDFQD1 \input_weight_reg[6][18]  ( .D(data_in[18]), .E(n429), .CP(clk), .Q(
        \input_weight[6][18] ) );
  EDFQD1 \input_weight_reg[6][17]  ( .D(data_in[17]), .E(n429), .CP(clk), .Q(
        \input_weight[6][17] ) );
  EDFQD1 \input_weight_reg[6][16]  ( .D(data_in[16]), .E(n429), .CP(clk), .Q(
        \input_weight[6][16] ) );
  EDFQD1 \input_weight_reg[6][15]  ( .D(data_in[15]), .E(n429), .CP(clk), .Q(
        \input_weight[6][15] ) );
  EDFQD1 \input_weight_reg[6][14]  ( .D(data_in[14]), .E(n429), .CP(clk), .Q(
        \input_weight[6][14] ) );
  EDFQD1 \input_weight_reg[6][13]  ( .D(data_in[13]), .E(n429), .CP(clk), .Q(
        \input_weight[6][13] ) );
  EDFQD1 \input_weight_reg[6][12]  ( .D(data_in[12]), .E(n428), .CP(clk), .Q(
        \input_weight[6][12] ) );
  EDFQD1 \input_weight_reg[6][11]  ( .D(data_in[11]), .E(n428), .CP(clk), .Q(
        \input_weight[6][11] ) );
  EDFQD1 \input_weight_reg[6][10]  ( .D(data_in[10]), .E(n428), .CP(clk), .Q(
        \input_weight[6][10] ) );
  EDFQD1 \input_weight_reg[6][9]  ( .D(data_in[9]), .E(n428), .CP(clk), .Q(
        \input_weight[6][9] ) );
  EDFQD1 \input_weight_reg[6][8]  ( .D(data_in[8]), .E(n428), .CP(clk), .Q(
        \input_weight[6][8] ) );
  EDFQD1 \input_weight_reg[6][7]  ( .D(data_in[7]), .E(n428), .CP(clk), .Q(
        \input_weight[6][7] ) );
  EDFQD1 \input_weight_reg[6][6]  ( .D(data_in[6]), .E(n428), .CP(clk), .Q(
        \input_weight[6][6] ) );
  EDFQD1 \input_weight_reg[6][5]  ( .D(data_in[5]), .E(n428), .CP(clk), .Q(
        \input_weight[6][5] ) );
  EDFQD1 \input_weight_reg[6][4]  ( .D(data_in[4]), .E(n428), .CP(clk), .Q(
        \input_weight[6][4] ) );
  EDFQD1 \input_weight_reg[6][3]  ( .D(data_in[3]), .E(n428), .CP(clk), .Q(
        \input_weight[6][3] ) );
  EDFQD1 \input_weight_reg[6][2]  ( .D(data_in[2]), .E(n428), .CP(clk), .Q(
        \input_weight[6][2] ) );
  EDFQD1 \input_weight_reg[6][1]  ( .D(data_in[1]), .E(n428), .CP(clk), .Q(
        \input_weight[6][1] ) );
  EDFQD1 \input_weight_reg[6][0]  ( .D(data_in[0]), .E(n428), .CP(clk), .Q(
        \input_weight[6][0] ) );
  EDFQD1 \input_value_reg[6][99]  ( .D(data_in[99]), .E(n317), .CP(clk), .Q(
        \input_value[6][99] ) );
  EDFQD1 \input_value_reg[6][100]  ( .D(data_in[100]), .E(n317), .CP(clk), .Q(
        \input_value[6][100] ) );
  EDFQD1 \input_value_reg[6][101]  ( .D(data_in[101]), .E(n317), .CP(clk), .Q(
        \input_value[6][101] ) );
  EDFQD1 \input_value_reg[6][102]  ( .D(data_in[102]), .E(n317), .CP(clk), .Q(
        \input_value[6][102] ) );
  EDFQD1 \input_value_reg[6][103]  ( .D(data_in[103]), .E(n317), .CP(clk), .Q(
        \input_value[6][103] ) );
  EDFQD1 \input_value_reg[6][104]  ( .D(data_in[104]), .E(n317), .CP(clk), .Q(
        \input_value[6][104] ) );
  EDFQD1 \input_value_reg[6][105]  ( .D(data_in[105]), .E(n317), .CP(clk), .Q(
        \input_value[6][105] ) );
  EDFQD1 \input_value_reg[6][106]  ( .D(data_in[106]), .E(n317), .CP(clk), .Q(
        \input_value[6][106] ) );
  EDFQD1 \input_value_reg[6][107]  ( .D(data_in[107]), .E(n317), .CP(clk), .Q(
        \input_value[6][107] ) );
  EDFQD1 \input_value_reg[6][108]  ( .D(data_in[108]), .E(n317), .CP(clk), .Q(
        \input_value[6][108] ) );
  EDFQD1 \input_value_reg[6][109]  ( .D(data_in[109]), .E(n317), .CP(clk), .Q(
        \input_value[6][109] ) );
  EDFQD1 \input_value_reg[6][110]  ( .D(data_in[110]), .E(n316), .CP(clk), .Q(
        \input_value[6][110] ) );
  EDFQD1 \input_value_reg[6][111]  ( .D(data_in[111]), .E(n316), .CP(clk), .Q(
        \input_value[6][111] ) );
  EDFQD1 \input_value_reg[6][112]  ( .D(data_in[112]), .E(n316), .CP(clk), .Q(
        \input_value[6][112] ) );
  EDFQD1 \input_value_reg[6][113]  ( .D(data_in[113]), .E(n316), .CP(clk), .Q(
        \input_value[6][113] ) );
  EDFQD1 \input_value_reg[6][114]  ( .D(data_in[114]), .E(n316), .CP(clk), .Q(
        \input_value[6][114] ) );
  EDFQD1 \input_value_reg[6][115]  ( .D(data_in[115]), .E(n316), .CP(clk), .Q(
        \input_value[6][115] ) );
  EDFQD1 \input_value_reg[6][116]  ( .D(data_in[116]), .E(n316), .CP(clk), .Q(
        \input_value[6][116] ) );
  EDFQD1 \input_value_reg[6][117]  ( .D(data_in[117]), .E(n316), .CP(clk), .Q(
        \input_value[6][117] ) );
  EDFQD1 \input_value_reg[6][118]  ( .D(data_in[118]), .E(n316), .CP(clk), .Q(
        \input_value[6][118] ) );
  EDFQD1 \input_value_reg[6][119]  ( .D(data_in[119]), .E(n316), .CP(clk), .Q(
        \input_value[6][119] ) );
  EDFQD1 \input_value_reg[6][120]  ( .D(data_in[120]), .E(n316), .CP(clk), .Q(
        \input_value[6][120] ) );
  EDFQD1 \input_value_reg[6][121]  ( .D(data_in[121]), .E(n316), .CP(clk), .Q(
        \input_value[6][121] ) );
  EDFQD1 \input_value_reg[6][122]  ( .D(data_in[122]), .E(n316), .CP(clk), .Q(
        \input_value[6][122] ) );
  EDFQD1 \input_value_reg[6][123]  ( .D(data_in[123]), .E(n315), .CP(clk), .Q(
        \input_value[6][123] ) );
  EDFQD1 \input_value_reg[6][124]  ( .D(data_in[124]), .E(n315), .CP(clk), .Q(
        \input_value[6][124] ) );
  EDFQD1 \input_value_reg[6][125]  ( .D(data_in[125]), .E(n315), .CP(clk), .Q(
        \input_value[6][125] ) );
  EDFQD1 \input_value_reg[6][126]  ( .D(data_in[126]), .E(n315), .CP(clk), .Q(
        \input_value[6][126] ) );
  EDFQD1 \input_value_reg[6][127]  ( .D(data_in[127]), .E(n315), .CP(clk), .Q(
        \input_value[6][127] ) );
  EDFQD1 \input_value_reg[6][98]  ( .D(data_in[98]), .E(n315), .CP(clk), .Q(
        \input_value[6][98] ) );
  EDFQD1 \input_value_reg[6][97]  ( .D(data_in[97]), .E(n315), .CP(clk), .Q(
        \input_value[6][97] ) );
  EDFQD1 \input_value_reg[6][96]  ( .D(data_in[96]), .E(n315), .CP(clk), .Q(
        \input_value[6][96] ) );
  EDFQD1 \input_value_reg[6][95]  ( .D(data_in[95]), .E(n315), .CP(clk), .Q(
        \input_value[6][95] ) );
  EDFQD1 \input_value_reg[6][94]  ( .D(data_in[94]), .E(n315), .CP(clk), .Q(
        \input_value[6][94] ) );
  EDFQD1 \input_value_reg[6][93]  ( .D(data_in[93]), .E(n315), .CP(clk), .Q(
        \input_value[6][93] ) );
  EDFQD1 \input_value_reg[6][92]  ( .D(data_in[92]), .E(n315), .CP(clk), .Q(
        \input_value[6][92] ) );
  EDFQD1 \input_value_reg[6][91]  ( .D(data_in[91]), .E(n315), .CP(clk), .Q(
        \input_value[6][91] ) );
  EDFQD1 \input_value_reg[6][90]  ( .D(data_in[90]), .E(n314), .CP(clk), .Q(
        \input_value[6][90] ) );
  EDFQD1 \input_value_reg[6][89]  ( .D(data_in[89]), .E(n314), .CP(clk), .Q(
        \input_value[6][89] ) );
  EDFQD1 \input_value_reg[6][88]  ( .D(data_in[88]), .E(n314), .CP(clk), .Q(
        \input_value[6][88] ) );
  EDFQD1 \input_value_reg[6][87]  ( .D(data_in[87]), .E(n314), .CP(clk), .Q(
        \input_value[6][87] ) );
  EDFQD1 \input_value_reg[6][86]  ( .D(data_in[86]), .E(n314), .CP(clk), .Q(
        \input_value[6][86] ) );
  EDFQD1 \input_value_reg[6][85]  ( .D(data_in[85]), .E(n314), .CP(clk), .Q(
        \input_value[6][85] ) );
  EDFQD1 \input_value_reg[6][84]  ( .D(data_in[84]), .E(n314), .CP(clk), .Q(
        \input_value[6][84] ) );
  EDFQD1 \input_value_reg[6][83]  ( .D(data_in[83]), .E(n314), .CP(clk), .Q(
        \input_value[6][83] ) );
  EDFQD1 \input_value_reg[6][82]  ( .D(data_in[82]), .E(n314), .CP(clk), .Q(
        \input_value[6][82] ) );
  EDFQD1 \input_value_reg[6][81]  ( .D(data_in[81]), .E(n314), .CP(clk), .Q(
        \input_value[6][81] ) );
  EDFQD1 \input_value_reg[6][80]  ( .D(data_in[80]), .E(n314), .CP(clk), .Q(
        \input_value[6][80] ) );
  EDFQD1 \input_value_reg[6][79]  ( .D(data_in[79]), .E(n314), .CP(clk), .Q(
        \input_value[6][79] ) );
  EDFQD1 \input_value_reg[6][78]  ( .D(data_in[78]), .E(n314), .CP(clk), .Q(
        \input_value[6][78] ) );
  EDFQD1 \input_value_reg[6][77]  ( .D(data_in[77]), .E(n313), .CP(clk), .Q(
        \input_value[6][77] ) );
  EDFQD1 \input_value_reg[6][76]  ( .D(data_in[76]), .E(n313), .CP(clk), .Q(
        \input_value[6][76] ) );
  EDFQD1 \input_value_reg[6][75]  ( .D(data_in[75]), .E(n313), .CP(clk), .Q(
        \input_value[6][75] ) );
  EDFQD1 \input_value_reg[6][74]  ( .D(data_in[74]), .E(n313), .CP(clk), .Q(
        \input_value[6][74] ) );
  EDFQD1 \input_value_reg[6][73]  ( .D(data_in[73]), .E(n313), .CP(clk), .Q(
        \input_value[6][73] ) );
  EDFQD1 \input_value_reg[6][72]  ( .D(data_in[72]), .E(n313), .CP(clk), .Q(
        \input_value[6][72] ) );
  EDFQD1 \input_value_reg[6][71]  ( .D(data_in[71]), .E(n313), .CP(clk), .Q(
        \input_value[6][71] ) );
  EDFQD1 \input_value_reg[6][70]  ( .D(data_in[70]), .E(n313), .CP(clk), .Q(
        \input_value[6][70] ) );
  EDFQD1 \input_value_reg[6][69]  ( .D(data_in[69]), .E(n313), .CP(clk), .Q(
        \input_value[6][69] ) );
  EDFQD1 \input_value_reg[6][68]  ( .D(data_in[68]), .E(n313), .CP(clk), .Q(
        \input_value[6][68] ) );
  EDFQD1 \input_value_reg[6][67]  ( .D(data_in[67]), .E(n313), .CP(clk), .Q(
        \input_value[6][67] ) );
  EDFQD1 \input_value_reg[6][66]  ( .D(data_in[66]), .E(n313), .CP(clk), .Q(
        \input_value[6][66] ) );
  EDFQD1 \input_value_reg[6][65]  ( .D(data_in[65]), .E(n313), .CP(clk), .Q(
        \input_value[6][65] ) );
  EDFQD1 \input_value_reg[6][64]  ( .D(data_in[64]), .E(n312), .CP(clk), .Q(
        \input_value[6][64] ) );
  EDFQD1 \input_value_reg[6][63]  ( .D(data_in[63]), .E(n312), .CP(clk), .Q(
        \input_value[6][63] ) );
  EDFQD1 \input_value_reg[6][62]  ( .D(data_in[62]), .E(n312), .CP(clk), .Q(
        \input_value[6][62] ) );
  EDFQD1 \input_value_reg[6][61]  ( .D(data_in[61]), .E(n312), .CP(clk), .Q(
        \input_value[6][61] ) );
  EDFQD1 \input_value_reg[6][60]  ( .D(data_in[60]), .E(n312), .CP(clk), .Q(
        \input_value[6][60] ) );
  EDFQD1 \input_value_reg[6][59]  ( .D(data_in[59]), .E(n312), .CP(clk), .Q(
        \input_value[6][59] ) );
  EDFQD1 \input_value_reg[6][58]  ( .D(data_in[58]), .E(n312), .CP(clk), .Q(
        \input_value[6][58] ) );
  EDFQD1 \input_value_reg[6][57]  ( .D(data_in[57]), .E(n312), .CP(clk), .Q(
        \input_value[6][57] ) );
  EDFQD1 \input_value_reg[6][56]  ( .D(data_in[56]), .E(n312), .CP(clk), .Q(
        \input_value[6][56] ) );
  EDFQD1 \input_value_reg[6][55]  ( .D(data_in[55]), .E(n312), .CP(clk), .Q(
        \input_value[6][55] ) );
  EDFQD1 \input_value_reg[6][54]  ( .D(data_in[54]), .E(n312), .CP(clk), .Q(
        \input_value[6][54] ) );
  EDFQD1 \input_value_reg[6][53]  ( .D(data_in[53]), .E(n312), .CP(clk), .Q(
        \input_value[6][53] ) );
  EDFQD1 \input_value_reg[6][52]  ( .D(data_in[52]), .E(n312), .CP(clk), .Q(
        \input_value[6][52] ) );
  EDFQD1 \input_value_reg[6][51]  ( .D(data_in[51]), .E(n311), .CP(clk), .Q(
        \input_value[6][51] ) );
  EDFQD1 \input_value_reg[6][50]  ( .D(data_in[50]), .E(n311), .CP(clk), .Q(
        \input_value[6][50] ) );
  EDFQD1 \input_value_reg[6][49]  ( .D(data_in[49]), .E(n311), .CP(clk), .Q(
        \input_value[6][49] ) );
  EDFQD1 \input_value_reg[6][48]  ( .D(data_in[48]), .E(n311), .CP(clk), .Q(
        \input_value[6][48] ) );
  EDFQD1 \input_value_reg[6][47]  ( .D(data_in[47]), .E(n311), .CP(clk), .Q(
        \input_value[6][47] ) );
  EDFQD1 \input_value_reg[6][46]  ( .D(data_in[46]), .E(n311), .CP(clk), .Q(
        \input_value[6][46] ) );
  EDFQD1 \input_value_reg[6][45]  ( .D(data_in[45]), .E(n311), .CP(clk), .Q(
        \input_value[6][45] ) );
  EDFQD1 \input_value_reg[6][44]  ( .D(data_in[44]), .E(n311), .CP(clk), .Q(
        \input_value[6][44] ) );
  EDFQD1 \input_value_reg[6][43]  ( .D(data_in[43]), .E(n311), .CP(clk), .Q(
        \input_value[6][43] ) );
  EDFQD1 \input_value_reg[6][42]  ( .D(data_in[42]), .E(n311), .CP(clk), .Q(
        \input_value[6][42] ) );
  EDFQD1 \input_value_reg[6][41]  ( .D(data_in[41]), .E(n311), .CP(clk), .Q(
        \input_value[6][41] ) );
  EDFQD1 \input_value_reg[6][40]  ( .D(data_in[40]), .E(n311), .CP(clk), .Q(
        \input_value[6][40] ) );
  EDFQD1 \input_value_reg[6][39]  ( .D(data_in[39]), .E(n311), .CP(clk), .Q(
        \input_value[6][39] ) );
  EDFQD1 \input_value_reg[6][38]  ( .D(data_in[38]), .E(n310), .CP(clk), .Q(
        \input_value[6][38] ) );
  EDFQD1 \input_value_reg[6][37]  ( .D(data_in[37]), .E(n310), .CP(clk), .Q(
        \input_value[6][37] ) );
  EDFQD1 \input_value_reg[6][36]  ( .D(data_in[36]), .E(n310), .CP(clk), .Q(
        \input_value[6][36] ) );
  EDFQD1 \input_value_reg[6][35]  ( .D(data_in[35]), .E(n310), .CP(clk), .Q(
        \input_value[6][35] ) );
  EDFQD1 \input_value_reg[6][34]  ( .D(data_in[34]), .E(n310), .CP(clk), .Q(
        \input_value[6][34] ) );
  EDFQD1 \input_value_reg[6][33]  ( .D(data_in[33]), .E(n310), .CP(clk), .Q(
        \input_value[6][33] ) );
  EDFQD1 \input_value_reg[6][32]  ( .D(data_in[32]), .E(n310), .CP(clk), .Q(
        \input_value[6][32] ) );
  EDFQD1 \input_value_reg[6][31]  ( .D(data_in[31]), .E(n310), .CP(clk), .Q(
        \input_value[6][31] ) );
  EDFQD1 \input_value_reg[6][30]  ( .D(data_in[30]), .E(n310), .CP(clk), .Q(
        \input_value[6][30] ) );
  EDFQD1 \input_value_reg[6][29]  ( .D(data_in[29]), .E(n310), .CP(clk), .Q(
        \input_value[6][29] ) );
  EDFQD1 \input_value_reg[6][28]  ( .D(data_in[28]), .E(n310), .CP(clk), .Q(
        \input_value[6][28] ) );
  EDFQD1 \input_value_reg[6][27]  ( .D(data_in[27]), .E(n310), .CP(clk), .Q(
        \input_value[6][27] ) );
  EDFQD1 \input_value_reg[6][26]  ( .D(data_in[26]), .E(n310), .CP(clk), .Q(
        \input_value[6][26] ) );
  EDFQD1 \input_value_reg[6][25]  ( .D(data_in[25]), .E(n309), .CP(clk), .Q(
        \input_value[6][25] ) );
  EDFQD1 \input_value_reg[6][24]  ( .D(data_in[24]), .E(n309), .CP(clk), .Q(
        \input_value[6][24] ) );
  EDFQD1 \input_value_reg[6][23]  ( .D(data_in[23]), .E(n309), .CP(clk), .Q(
        \input_value[6][23] ) );
  EDFQD1 \input_value_reg[6][22]  ( .D(data_in[22]), .E(n309), .CP(clk), .Q(
        \input_value[6][22] ) );
  EDFQD1 \input_value_reg[6][21]  ( .D(data_in[21]), .E(n309), .CP(clk), .Q(
        \input_value[6][21] ) );
  EDFQD1 \input_value_reg[6][20]  ( .D(data_in[20]), .E(n309), .CP(clk), .Q(
        \input_value[6][20] ) );
  EDFQD1 \input_value_reg[6][19]  ( .D(data_in[19]), .E(n309), .CP(clk), .Q(
        \input_value[6][19] ) );
  EDFQD1 \input_value_reg[6][18]  ( .D(data_in[18]), .E(n309), .CP(clk), .Q(
        \input_value[6][18] ) );
  EDFQD1 \input_value_reg[6][17]  ( .D(data_in[17]), .E(n309), .CP(clk), .Q(
        \input_value[6][17] ) );
  EDFQD1 \input_value_reg[6][16]  ( .D(data_in[16]), .E(n309), .CP(clk), .Q(
        \input_value[6][16] ) );
  EDFQD1 \input_value_reg[6][15]  ( .D(data_in[15]), .E(n309), .CP(clk), .Q(
        \input_value[6][15] ) );
  EDFQD1 \input_value_reg[6][14]  ( .D(data_in[14]), .E(n309), .CP(clk), .Q(
        \input_value[6][14] ) );
  EDFQD1 \input_value_reg[6][13]  ( .D(data_in[13]), .E(n309), .CP(clk), .Q(
        \input_value[6][13] ) );
  EDFQD1 \input_value_reg[6][12]  ( .D(data_in[12]), .E(n308), .CP(clk), .Q(
        \input_value[6][12] ) );
  EDFQD1 \input_value_reg[6][11]  ( .D(data_in[11]), .E(n308), .CP(clk), .Q(
        \input_value[6][11] ) );
  EDFQD1 \input_value_reg[6][10]  ( .D(data_in[10]), .E(n308), .CP(clk), .Q(
        \input_value[6][10] ) );
  EDFQD1 \input_value_reg[6][9]  ( .D(data_in[9]), .E(n308), .CP(clk), .Q(
        \input_value[6][9] ) );
  EDFQD1 \input_value_reg[6][8]  ( .D(data_in[8]), .E(n308), .CP(clk), .Q(
        \input_value[6][8] ) );
  EDFQD1 \input_value_reg[6][7]  ( .D(data_in[7]), .E(n308), .CP(clk), .Q(
        \input_value[6][7] ) );
  EDFQD1 \input_value_reg[6][6]  ( .D(data_in[6]), .E(n308), .CP(clk), .Q(
        \input_value[6][6] ) );
  EDFQD1 \input_value_reg[6][5]  ( .D(data_in[5]), .E(n308), .CP(clk), .Q(
        \input_value[6][5] ) );
  EDFQD1 \input_value_reg[6][4]  ( .D(data_in[4]), .E(n308), .CP(clk), .Q(
        \input_value[6][4] ) );
  EDFQD1 \input_value_reg[6][3]  ( .D(data_in[3]), .E(n308), .CP(clk), .Q(
        \input_value[6][3] ) );
  EDFQD1 \input_value_reg[6][2]  ( .D(data_in[2]), .E(n308), .CP(clk), .Q(
        \input_value[6][2] ) );
  EDFQD1 \input_value_reg[6][1]  ( .D(data_in[1]), .E(n308), .CP(clk), .Q(
        \input_value[6][1] ) );
  EDFQD1 \input_value_reg[6][0]  ( .D(data_in[0]), .E(n308), .CP(clk), .Q(
        \input_value[6][0] ) );
  EDFQD1 \input_value_reg[2][99]  ( .D(data_in[99]), .E(n377), .CP(clk), .Q(
        \input_value[2][99] ) );
  EDFQD1 \input_value_reg[2][100]  ( .D(data_in[100]), .E(n377), .CP(clk), .Q(
        \input_value[2][100] ) );
  EDFQD1 \input_value_reg[2][101]  ( .D(data_in[101]), .E(n377), .CP(clk), .Q(
        \input_value[2][101] ) );
  EDFQD1 \input_value_reg[2][102]  ( .D(data_in[102]), .E(n377), .CP(clk), .Q(
        \input_value[2][102] ) );
  EDFQD1 \input_value_reg[2][103]  ( .D(data_in[103]), .E(n377), .CP(clk), .Q(
        \input_value[2][103] ) );
  EDFQD1 \input_value_reg[2][104]  ( .D(data_in[104]), .E(n377), .CP(clk), .Q(
        \input_value[2][104] ) );
  EDFQD1 \input_value_reg[2][105]  ( .D(data_in[105]), .E(n377), .CP(clk), .Q(
        \input_value[2][105] ) );
  EDFQD1 \input_value_reg[2][106]  ( .D(data_in[106]), .E(n377), .CP(clk), .Q(
        \input_value[2][106] ) );
  EDFQD1 \input_value_reg[2][107]  ( .D(data_in[107]), .E(n377), .CP(clk), .Q(
        \input_value[2][107] ) );
  EDFQD1 \input_value_reg[2][108]  ( .D(data_in[108]), .E(n377), .CP(clk), .Q(
        \input_value[2][108] ) );
  EDFQD1 \input_value_reg[2][109]  ( .D(data_in[109]), .E(n377), .CP(clk), .Q(
        \input_value[2][109] ) );
  EDFQD1 \input_value_reg[2][110]  ( .D(data_in[110]), .E(n376), .CP(clk), .Q(
        \input_value[2][110] ) );
  EDFQD1 \input_value_reg[2][111]  ( .D(data_in[111]), .E(n376), .CP(clk), .Q(
        \input_value[2][111] ) );
  EDFQD1 \input_value_reg[2][112]  ( .D(data_in[112]), .E(n376), .CP(clk), .Q(
        \input_value[2][112] ) );
  EDFQD1 \input_value_reg[2][113]  ( .D(data_in[113]), .E(n376), .CP(clk), .Q(
        \input_value[2][113] ) );
  EDFQD1 \input_value_reg[2][114]  ( .D(data_in[114]), .E(n376), .CP(clk), .Q(
        \input_value[2][114] ) );
  EDFQD1 \input_value_reg[2][115]  ( .D(data_in[115]), .E(n376), .CP(clk), .Q(
        \input_value[2][115] ) );
  EDFQD1 \input_value_reg[2][116]  ( .D(data_in[116]), .E(n376), .CP(clk), .Q(
        \input_value[2][116] ) );
  EDFQD1 \input_value_reg[2][117]  ( .D(data_in[117]), .E(n376), .CP(clk), .Q(
        \input_value[2][117] ) );
  EDFQD1 \input_value_reg[2][118]  ( .D(data_in[118]), .E(n376), .CP(clk), .Q(
        \input_value[2][118] ) );
  EDFQD1 \input_value_reg[2][119]  ( .D(data_in[119]), .E(n376), .CP(clk), .Q(
        \input_value[2][119] ) );
  EDFQD1 \input_value_reg[2][120]  ( .D(data_in[120]), .E(n376), .CP(clk), .Q(
        \input_value[2][120] ) );
  EDFQD1 \input_value_reg[2][121]  ( .D(data_in[121]), .E(n376), .CP(clk), .Q(
        \input_value[2][121] ) );
  EDFQD1 \input_value_reg[2][122]  ( .D(data_in[122]), .E(n376), .CP(clk), .Q(
        \input_value[2][122] ) );
  EDFQD1 \input_value_reg[2][123]  ( .D(data_in[123]), .E(n375), .CP(clk), .Q(
        \input_value[2][123] ) );
  EDFQD1 \input_value_reg[2][124]  ( .D(data_in[124]), .E(n375), .CP(clk), .Q(
        \input_value[2][124] ) );
  EDFQD1 \input_value_reg[2][125]  ( .D(data_in[125]), .E(n375), .CP(clk), .Q(
        \input_value[2][125] ) );
  EDFQD1 \input_value_reg[2][126]  ( .D(data_in[126]), .E(n375), .CP(clk), .Q(
        \input_value[2][126] ) );
  EDFQD1 \input_value_reg[2][127]  ( .D(data_in[127]), .E(n375), .CP(clk), .Q(
        \input_value[2][127] ) );
  EDFQD1 \input_value_reg[2][98]  ( .D(data_in[98]), .E(n375), .CP(clk), .Q(
        \input_value[2][98] ) );
  EDFQD1 \input_value_reg[2][97]  ( .D(data_in[97]), .E(n375), .CP(clk), .Q(
        \input_value[2][97] ) );
  EDFQD1 \input_value_reg[2][96]  ( .D(data_in[96]), .E(n375), .CP(clk), .Q(
        \input_value[2][96] ) );
  EDFQD1 \input_value_reg[2][95]  ( .D(data_in[95]), .E(n375), .CP(clk), .Q(
        \input_value[2][95] ) );
  EDFQD1 \input_value_reg[2][94]  ( .D(data_in[94]), .E(n375), .CP(clk), .Q(
        \input_value[2][94] ) );
  EDFQD1 \input_value_reg[2][93]  ( .D(data_in[93]), .E(n375), .CP(clk), .Q(
        \input_value[2][93] ) );
  EDFQD1 \input_value_reg[2][92]  ( .D(data_in[92]), .E(n375), .CP(clk), .Q(
        \input_value[2][92] ) );
  EDFQD1 \input_value_reg[2][91]  ( .D(data_in[91]), .E(n375), .CP(clk), .Q(
        \input_value[2][91] ) );
  EDFQD1 \input_value_reg[2][90]  ( .D(data_in[90]), .E(n374), .CP(clk), .Q(
        \input_value[2][90] ) );
  EDFQD1 \input_value_reg[2][89]  ( .D(data_in[89]), .E(n374), .CP(clk), .Q(
        \input_value[2][89] ) );
  EDFQD1 \input_value_reg[2][88]  ( .D(data_in[88]), .E(n374), .CP(clk), .Q(
        \input_value[2][88] ) );
  EDFQD1 \input_value_reg[2][87]  ( .D(data_in[87]), .E(n374), .CP(clk), .Q(
        \input_value[2][87] ) );
  EDFQD1 \input_value_reg[2][86]  ( .D(data_in[86]), .E(n374), .CP(clk), .Q(
        \input_value[2][86] ) );
  EDFQD1 \input_value_reg[2][85]  ( .D(data_in[85]), .E(n374), .CP(clk), .Q(
        \input_value[2][85] ) );
  EDFQD1 \input_value_reg[2][84]  ( .D(data_in[84]), .E(n374), .CP(clk), .Q(
        \input_value[2][84] ) );
  EDFQD1 \input_value_reg[2][83]  ( .D(data_in[83]), .E(n374), .CP(clk), .Q(
        \input_value[2][83] ) );
  EDFQD1 \input_value_reg[2][82]  ( .D(data_in[82]), .E(n374), .CP(clk), .Q(
        \input_value[2][82] ) );
  EDFQD1 \input_value_reg[2][81]  ( .D(data_in[81]), .E(n374), .CP(clk), .Q(
        \input_value[2][81] ) );
  EDFQD1 \input_value_reg[2][80]  ( .D(data_in[80]), .E(n374), .CP(clk), .Q(
        \input_value[2][80] ) );
  EDFQD1 \input_value_reg[2][79]  ( .D(data_in[79]), .E(n374), .CP(clk), .Q(
        \input_value[2][79] ) );
  EDFQD1 \input_value_reg[2][78]  ( .D(data_in[78]), .E(n374), .CP(clk), .Q(
        \input_value[2][78] ) );
  EDFQD1 \input_value_reg[2][77]  ( .D(data_in[77]), .E(n373), .CP(clk), .Q(
        \input_value[2][77] ) );
  EDFQD1 \input_value_reg[2][76]  ( .D(data_in[76]), .E(n373), .CP(clk), .Q(
        \input_value[2][76] ) );
  EDFQD1 \input_value_reg[2][75]  ( .D(data_in[75]), .E(n373), .CP(clk), .Q(
        \input_value[2][75] ) );
  EDFQD1 \input_value_reg[2][74]  ( .D(data_in[74]), .E(n373), .CP(clk), .Q(
        \input_value[2][74] ) );
  EDFQD1 \input_value_reg[2][73]  ( .D(data_in[73]), .E(n373), .CP(clk), .Q(
        \input_value[2][73] ) );
  EDFQD1 \input_value_reg[2][72]  ( .D(data_in[72]), .E(n373), .CP(clk), .Q(
        \input_value[2][72] ) );
  EDFQD1 \input_value_reg[2][71]  ( .D(data_in[71]), .E(n373), .CP(clk), .Q(
        \input_value[2][71] ) );
  EDFQD1 \input_value_reg[2][70]  ( .D(data_in[70]), .E(n373), .CP(clk), .Q(
        \input_value[2][70] ) );
  EDFQD1 \input_value_reg[2][69]  ( .D(data_in[69]), .E(n373), .CP(clk), .Q(
        \input_value[2][69] ) );
  EDFQD1 \input_value_reg[2][68]  ( .D(data_in[68]), .E(n373), .CP(clk), .Q(
        \input_value[2][68] ) );
  EDFQD1 \input_value_reg[2][67]  ( .D(data_in[67]), .E(n373), .CP(clk), .Q(
        \input_value[2][67] ) );
  EDFQD1 \input_value_reg[2][66]  ( .D(data_in[66]), .E(n373), .CP(clk), .Q(
        \input_value[2][66] ) );
  EDFQD1 \input_value_reg[2][65]  ( .D(data_in[65]), .E(n373), .CP(clk), .Q(
        \input_value[2][65] ) );
  EDFQD1 \input_value_reg[2][64]  ( .D(data_in[64]), .E(n372), .CP(clk), .Q(
        \input_value[2][64] ) );
  EDFQD1 \input_value_reg[2][63]  ( .D(data_in[63]), .E(n372), .CP(clk), .Q(
        \input_value[2][63] ) );
  EDFQD1 \input_value_reg[2][62]  ( .D(data_in[62]), .E(n372), .CP(clk), .Q(
        \input_value[2][62] ) );
  EDFQD1 \input_value_reg[2][61]  ( .D(data_in[61]), .E(n372), .CP(clk), .Q(
        \input_value[2][61] ) );
  EDFQD1 \input_value_reg[2][60]  ( .D(data_in[60]), .E(n372), .CP(clk), .Q(
        \input_value[2][60] ) );
  EDFQD1 \input_value_reg[2][59]  ( .D(data_in[59]), .E(n372), .CP(clk), .Q(
        \input_value[2][59] ) );
  EDFQD1 \input_value_reg[2][58]  ( .D(data_in[58]), .E(n372), .CP(clk), .Q(
        \input_value[2][58] ) );
  EDFQD1 \input_value_reg[2][57]  ( .D(data_in[57]), .E(n372), .CP(clk), .Q(
        \input_value[2][57] ) );
  EDFQD1 \input_value_reg[2][56]  ( .D(data_in[56]), .E(n372), .CP(clk), .Q(
        \input_value[2][56] ) );
  EDFQD1 \input_value_reg[2][55]  ( .D(data_in[55]), .E(n372), .CP(clk), .Q(
        \input_value[2][55] ) );
  EDFQD1 \input_value_reg[2][54]  ( .D(data_in[54]), .E(n372), .CP(clk), .Q(
        \input_value[2][54] ) );
  EDFQD1 \input_value_reg[2][53]  ( .D(data_in[53]), .E(n372), .CP(clk), .Q(
        \input_value[2][53] ) );
  EDFQD1 \input_value_reg[2][52]  ( .D(data_in[52]), .E(n372), .CP(clk), .Q(
        \input_value[2][52] ) );
  EDFQD1 \input_value_reg[2][51]  ( .D(data_in[51]), .E(n371), .CP(clk), .Q(
        \input_value[2][51] ) );
  EDFQD1 \input_value_reg[2][50]  ( .D(data_in[50]), .E(n371), .CP(clk), .Q(
        \input_value[2][50] ) );
  EDFQD1 \input_value_reg[2][49]  ( .D(data_in[49]), .E(n371), .CP(clk), .Q(
        \input_value[2][49] ) );
  EDFQD1 \input_value_reg[2][48]  ( .D(data_in[48]), .E(n371), .CP(clk), .Q(
        \input_value[2][48] ) );
  EDFQD1 \input_value_reg[2][47]  ( .D(data_in[47]), .E(n371), .CP(clk), .Q(
        \input_value[2][47] ) );
  EDFQD1 \input_value_reg[2][46]  ( .D(data_in[46]), .E(n371), .CP(clk), .Q(
        \input_value[2][46] ) );
  EDFQD1 \input_value_reg[2][45]  ( .D(data_in[45]), .E(n371), .CP(clk), .Q(
        \input_value[2][45] ) );
  EDFQD1 \input_value_reg[2][44]  ( .D(data_in[44]), .E(n371), .CP(clk), .Q(
        \input_value[2][44] ) );
  EDFQD1 \input_value_reg[2][43]  ( .D(data_in[43]), .E(n371), .CP(clk), .Q(
        \input_value[2][43] ) );
  EDFQD1 \input_value_reg[2][42]  ( .D(data_in[42]), .E(n371), .CP(clk), .Q(
        \input_value[2][42] ) );
  EDFQD1 \input_value_reg[2][41]  ( .D(data_in[41]), .E(n371), .CP(clk), .Q(
        \input_value[2][41] ) );
  EDFQD1 \input_value_reg[2][40]  ( .D(data_in[40]), .E(n371), .CP(clk), .Q(
        \input_value[2][40] ) );
  EDFQD1 \input_value_reg[2][39]  ( .D(data_in[39]), .E(n371), .CP(clk), .Q(
        \input_value[2][39] ) );
  EDFQD1 \input_value_reg[2][38]  ( .D(data_in[38]), .E(n370), .CP(clk), .Q(
        \input_value[2][38] ) );
  EDFQD1 \input_value_reg[2][37]  ( .D(data_in[37]), .E(n370), .CP(clk), .Q(
        \input_value[2][37] ) );
  EDFQD1 \input_value_reg[2][36]  ( .D(data_in[36]), .E(n370), .CP(clk), .Q(
        \input_value[2][36] ) );
  EDFQD1 \input_value_reg[2][35]  ( .D(data_in[35]), .E(n370), .CP(clk), .Q(
        \input_value[2][35] ) );
  EDFQD1 \input_value_reg[2][34]  ( .D(data_in[34]), .E(n370), .CP(clk), .Q(
        \input_value[2][34] ) );
  EDFQD1 \input_value_reg[2][33]  ( .D(data_in[33]), .E(n370), .CP(clk), .Q(
        \input_value[2][33] ) );
  EDFQD1 \input_value_reg[2][32]  ( .D(data_in[32]), .E(n370), .CP(clk), .Q(
        \input_value[2][32] ) );
  EDFQD1 \input_value_reg[2][31]  ( .D(data_in[31]), .E(n370), .CP(clk), .Q(
        \input_value[2][31] ) );
  EDFQD1 \input_value_reg[2][30]  ( .D(data_in[30]), .E(n370), .CP(clk), .Q(
        \input_value[2][30] ) );
  EDFQD1 \input_value_reg[2][29]  ( .D(data_in[29]), .E(n370), .CP(clk), .Q(
        \input_value[2][29] ) );
  EDFQD1 \input_value_reg[2][28]  ( .D(data_in[28]), .E(n370), .CP(clk), .Q(
        \input_value[2][28] ) );
  EDFQD1 \input_value_reg[2][27]  ( .D(data_in[27]), .E(n370), .CP(clk), .Q(
        \input_value[2][27] ) );
  EDFQD1 \input_value_reg[2][26]  ( .D(data_in[26]), .E(n370), .CP(clk), .Q(
        \input_value[2][26] ) );
  EDFQD1 \input_value_reg[2][25]  ( .D(data_in[25]), .E(n369), .CP(clk), .Q(
        \input_value[2][25] ) );
  EDFQD1 \input_value_reg[2][24]  ( .D(data_in[24]), .E(n369), .CP(clk), .Q(
        \input_value[2][24] ) );
  EDFQD1 \input_value_reg[2][23]  ( .D(data_in[23]), .E(n369), .CP(clk), .Q(
        \input_value[2][23] ) );
  EDFQD1 \input_value_reg[2][22]  ( .D(data_in[22]), .E(n369), .CP(clk), .Q(
        \input_value[2][22] ) );
  EDFQD1 \input_value_reg[2][21]  ( .D(data_in[21]), .E(n369), .CP(clk), .Q(
        \input_value[2][21] ) );
  EDFQD1 \input_value_reg[2][20]  ( .D(data_in[20]), .E(n369), .CP(clk), .Q(
        \input_value[2][20] ) );
  EDFQD1 \input_value_reg[2][19]  ( .D(data_in[19]), .E(n369), .CP(clk), .Q(
        \input_value[2][19] ) );
  EDFQD1 \input_value_reg[2][18]  ( .D(data_in[18]), .E(n369), .CP(clk), .Q(
        \input_value[2][18] ) );
  EDFQD1 \input_value_reg[2][17]  ( .D(data_in[17]), .E(n369), .CP(clk), .Q(
        \input_value[2][17] ) );
  EDFQD1 \input_value_reg[2][16]  ( .D(data_in[16]), .E(n369), .CP(clk), .Q(
        \input_value[2][16] ) );
  EDFQD1 \input_value_reg[2][15]  ( .D(data_in[15]), .E(n369), .CP(clk), .Q(
        \input_value[2][15] ) );
  EDFQD1 \input_value_reg[2][14]  ( .D(data_in[14]), .E(n369), .CP(clk), .Q(
        \input_value[2][14] ) );
  EDFQD1 \input_value_reg[2][13]  ( .D(data_in[13]), .E(n369), .CP(clk), .Q(
        \input_value[2][13] ) );
  EDFQD1 \input_value_reg[2][12]  ( .D(data_in[12]), .E(n368), .CP(clk), .Q(
        \input_value[2][12] ) );
  EDFQD1 \input_value_reg[2][11]  ( .D(data_in[11]), .E(n368), .CP(clk), .Q(
        \input_value[2][11] ) );
  EDFQD1 \input_value_reg[2][10]  ( .D(data_in[10]), .E(n368), .CP(clk), .Q(
        \input_value[2][10] ) );
  EDFQD1 \input_value_reg[2][9]  ( .D(data_in[9]), .E(n368), .CP(clk), .Q(
        \input_value[2][9] ) );
  EDFQD1 \input_value_reg[2][8]  ( .D(data_in[8]), .E(n368), .CP(clk), .Q(
        \input_value[2][8] ) );
  EDFQD1 \input_value_reg[2][7]  ( .D(data_in[7]), .E(n368), .CP(clk), .Q(
        \input_value[2][7] ) );
  EDFQD1 \input_value_reg[2][6]  ( .D(data_in[6]), .E(n368), .CP(clk), .Q(
        \input_value[2][6] ) );
  EDFQD1 \input_value_reg[2][5]  ( .D(data_in[5]), .E(n368), .CP(clk), .Q(
        \input_value[2][5] ) );
  EDFQD1 \input_value_reg[2][4]  ( .D(data_in[4]), .E(n368), .CP(clk), .Q(
        \input_value[2][4] ) );
  EDFQD1 \input_value_reg[2][3]  ( .D(data_in[3]), .E(n368), .CP(clk), .Q(
        \input_value[2][3] ) );
  EDFQD1 \input_value_reg[2][2]  ( .D(data_in[2]), .E(n368), .CP(clk), .Q(
        \input_value[2][2] ) );
  EDFQD1 \input_value_reg[2][1]  ( .D(data_in[1]), .E(n368), .CP(clk), .Q(
        \input_value[2][1] ) );
  EDFQD1 \input_value_reg[2][0]  ( .D(data_in[0]), .E(n368), .CP(clk), .Q(
        \input_value[2][0] ) );
  EDFQD1 \input_weight_reg[2][99]  ( .D(data_in[99]), .E(n497), .CP(clk), .Q(
        \input_weight[2][99] ) );
  EDFQD1 \input_weight_reg[2][100]  ( .D(data_in[100]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][100] ) );
  EDFQD1 \input_weight_reg[2][101]  ( .D(data_in[101]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][101] ) );
  EDFQD1 \input_weight_reg[2][102]  ( .D(data_in[102]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][102] ) );
  EDFQD1 \input_weight_reg[2][103]  ( .D(data_in[103]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][103] ) );
  EDFQD1 \input_weight_reg[2][104]  ( .D(data_in[104]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][104] ) );
  EDFQD1 \input_weight_reg[2][105]  ( .D(data_in[105]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][105] ) );
  EDFQD1 \input_weight_reg[2][106]  ( .D(data_in[106]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][106] ) );
  EDFQD1 \input_weight_reg[2][107]  ( .D(data_in[107]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][107] ) );
  EDFQD1 \input_weight_reg[2][108]  ( .D(data_in[108]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][108] ) );
  EDFQD1 \input_weight_reg[2][109]  ( .D(data_in[109]), .E(n497), .CP(clk), 
        .Q(\input_weight[2][109] ) );
  EDFQD1 \input_weight_reg[2][110]  ( .D(data_in[110]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][110] ) );
  EDFQD1 \input_weight_reg[2][111]  ( .D(data_in[111]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][111] ) );
  EDFQD1 \input_weight_reg[2][112]  ( .D(data_in[112]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][112] ) );
  EDFQD1 \input_weight_reg[2][113]  ( .D(data_in[113]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][113] ) );
  EDFQD1 \input_weight_reg[2][114]  ( .D(data_in[114]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][114] ) );
  EDFQD1 \input_weight_reg[2][115]  ( .D(data_in[115]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][115] ) );
  EDFQD1 \input_weight_reg[2][116]  ( .D(data_in[116]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][116] ) );
  EDFQD1 \input_weight_reg[2][117]  ( .D(data_in[117]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][117] ) );
  EDFQD1 \input_weight_reg[2][118]  ( .D(data_in[118]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][118] ) );
  EDFQD1 \input_weight_reg[2][119]  ( .D(data_in[119]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][119] ) );
  EDFQD1 \input_weight_reg[2][120]  ( .D(data_in[120]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][120] ) );
  EDFQD1 \input_weight_reg[2][121]  ( .D(data_in[121]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][121] ) );
  EDFQD1 \input_weight_reg[2][122]  ( .D(data_in[122]), .E(n496), .CP(clk), 
        .Q(\input_weight[2][122] ) );
  EDFQD1 \input_weight_reg[2][123]  ( .D(data_in[123]), .E(n495), .CP(clk), 
        .Q(\input_weight[2][123] ) );
  EDFQD1 \input_weight_reg[2][124]  ( .D(data_in[124]), .E(n495), .CP(clk), 
        .Q(\input_weight[2][124] ) );
  EDFQD1 \input_weight_reg[2][125]  ( .D(data_in[125]), .E(n495), .CP(clk), 
        .Q(\input_weight[2][125] ) );
  EDFQD1 \input_weight_reg[2][126]  ( .D(data_in[126]), .E(n495), .CP(clk), 
        .Q(\input_weight[2][126] ) );
  EDFQD1 \input_weight_reg[2][127]  ( .D(data_in[127]), .E(n495), .CP(clk), 
        .Q(\input_weight[2][127] ) );
  EDFQD1 \input_weight_reg[2][98]  ( .D(data_in[98]), .E(n495), .CP(clk), .Q(
        \input_weight[2][98] ) );
  EDFQD1 \input_weight_reg[2][97]  ( .D(data_in[97]), .E(n495), .CP(clk), .Q(
        \input_weight[2][97] ) );
  EDFQD1 \input_weight_reg[2][96]  ( .D(data_in[96]), .E(n495), .CP(clk), .Q(
        \input_weight[2][96] ) );
  EDFQD1 \input_weight_reg[2][95]  ( .D(data_in[95]), .E(n495), .CP(clk), .Q(
        \input_weight[2][95] ) );
  EDFQD1 \input_weight_reg[2][94]  ( .D(data_in[94]), .E(n495), .CP(clk), .Q(
        \input_weight[2][94] ) );
  EDFQD1 \input_weight_reg[2][93]  ( .D(data_in[93]), .E(n495), .CP(clk), .Q(
        \input_weight[2][93] ) );
  EDFQD1 \input_weight_reg[2][92]  ( .D(data_in[92]), .E(n495), .CP(clk), .Q(
        \input_weight[2][92] ) );
  EDFQD1 \input_weight_reg[2][91]  ( .D(data_in[91]), .E(n495), .CP(clk), .Q(
        \input_weight[2][91] ) );
  EDFQD1 \input_weight_reg[2][90]  ( .D(data_in[90]), .E(n494), .CP(clk), .Q(
        \input_weight[2][90] ) );
  EDFQD1 \input_weight_reg[2][89]  ( .D(data_in[89]), .E(n494), .CP(clk), .Q(
        \input_weight[2][89] ) );
  EDFQD1 \input_weight_reg[2][88]  ( .D(data_in[88]), .E(n494), .CP(clk), .Q(
        \input_weight[2][88] ) );
  EDFQD1 \input_weight_reg[2][87]  ( .D(data_in[87]), .E(n494), .CP(clk), .Q(
        \input_weight[2][87] ) );
  EDFQD1 \input_weight_reg[2][86]  ( .D(data_in[86]), .E(n494), .CP(clk), .Q(
        \input_weight[2][86] ) );
  EDFQD1 \input_weight_reg[2][85]  ( .D(data_in[85]), .E(n494), .CP(clk), .Q(
        \input_weight[2][85] ) );
  EDFQD1 \input_weight_reg[2][84]  ( .D(data_in[84]), .E(n494), .CP(clk), .Q(
        \input_weight[2][84] ) );
  EDFQD1 \input_weight_reg[2][83]  ( .D(data_in[83]), .E(n494), .CP(clk), .Q(
        \input_weight[2][83] ) );
  EDFQD1 \input_weight_reg[2][82]  ( .D(data_in[82]), .E(n494), .CP(clk), .Q(
        \input_weight[2][82] ) );
  EDFQD1 \input_weight_reg[2][81]  ( .D(data_in[81]), .E(n494), .CP(clk), .Q(
        \input_weight[2][81] ) );
  EDFQD1 \input_weight_reg[2][80]  ( .D(data_in[80]), .E(n494), .CP(clk), .Q(
        \input_weight[2][80] ) );
  EDFQD1 \input_weight_reg[2][79]  ( .D(data_in[79]), .E(n494), .CP(clk), .Q(
        \input_weight[2][79] ) );
  EDFQD1 \input_weight_reg[2][78]  ( .D(data_in[78]), .E(n494), .CP(clk), .Q(
        \input_weight[2][78] ) );
  EDFQD1 \input_weight_reg[2][77]  ( .D(data_in[77]), .E(n493), .CP(clk), .Q(
        \input_weight[2][77] ) );
  EDFQD1 \input_weight_reg[2][76]  ( .D(data_in[76]), .E(n493), .CP(clk), .Q(
        \input_weight[2][76] ) );
  EDFQD1 \input_weight_reg[2][75]  ( .D(data_in[75]), .E(n493), .CP(clk), .Q(
        \input_weight[2][75] ) );
  EDFQD1 \input_weight_reg[2][74]  ( .D(data_in[74]), .E(n493), .CP(clk), .Q(
        \input_weight[2][74] ) );
  EDFQD1 \input_weight_reg[2][73]  ( .D(data_in[73]), .E(n493), .CP(clk), .Q(
        \input_weight[2][73] ) );
  EDFQD1 \input_weight_reg[2][72]  ( .D(data_in[72]), .E(n493), .CP(clk), .Q(
        \input_weight[2][72] ) );
  EDFQD1 \input_weight_reg[2][71]  ( .D(data_in[71]), .E(n493), .CP(clk), .Q(
        \input_weight[2][71] ) );
  EDFQD1 \input_weight_reg[2][70]  ( .D(data_in[70]), .E(n493), .CP(clk), .Q(
        \input_weight[2][70] ) );
  EDFQD1 \input_weight_reg[2][69]  ( .D(data_in[69]), .E(n493), .CP(clk), .Q(
        \input_weight[2][69] ) );
  EDFQD1 \input_weight_reg[2][68]  ( .D(data_in[68]), .E(n493), .CP(clk), .Q(
        \input_weight[2][68] ) );
  EDFQD1 \input_weight_reg[2][67]  ( .D(data_in[67]), .E(n493), .CP(clk), .Q(
        \input_weight[2][67] ) );
  EDFQD1 \input_weight_reg[2][66]  ( .D(data_in[66]), .E(n493), .CP(clk), .Q(
        \input_weight[2][66] ) );
  EDFQD1 \input_weight_reg[2][65]  ( .D(data_in[65]), .E(n493), .CP(clk), .Q(
        \input_weight[2][65] ) );
  EDFQD1 \input_weight_reg[2][64]  ( .D(data_in[64]), .E(n492), .CP(clk), .Q(
        \input_weight[2][64] ) );
  EDFQD1 \input_weight_reg[2][63]  ( .D(data_in[63]), .E(n492), .CP(clk), .Q(
        \input_weight[2][63] ) );
  EDFQD1 \input_weight_reg[2][62]  ( .D(data_in[62]), .E(n492), .CP(clk), .Q(
        \input_weight[2][62] ) );
  EDFQD1 \input_weight_reg[2][61]  ( .D(data_in[61]), .E(n492), .CP(clk), .Q(
        \input_weight[2][61] ) );
  EDFQD1 \input_weight_reg[2][60]  ( .D(data_in[60]), .E(n492), .CP(clk), .Q(
        \input_weight[2][60] ) );
  EDFQD1 \input_weight_reg[2][59]  ( .D(data_in[59]), .E(n492), .CP(clk), .Q(
        \input_weight[2][59] ) );
  EDFQD1 \input_weight_reg[2][58]  ( .D(data_in[58]), .E(n492), .CP(clk), .Q(
        \input_weight[2][58] ) );
  EDFQD1 \input_weight_reg[2][57]  ( .D(data_in[57]), .E(n492), .CP(clk), .Q(
        \input_weight[2][57] ) );
  EDFQD1 \input_weight_reg[2][56]  ( .D(data_in[56]), .E(n492), .CP(clk), .Q(
        \input_weight[2][56] ) );
  EDFQD1 \input_weight_reg[2][55]  ( .D(data_in[55]), .E(n492), .CP(clk), .Q(
        \input_weight[2][55] ) );
  EDFQD1 \input_weight_reg[2][54]  ( .D(data_in[54]), .E(n492), .CP(clk), .Q(
        \input_weight[2][54] ) );
  EDFQD1 \input_weight_reg[2][53]  ( .D(data_in[53]), .E(n492), .CP(clk), .Q(
        \input_weight[2][53] ) );
  EDFQD1 \input_weight_reg[2][52]  ( .D(data_in[52]), .E(n492), .CP(clk), .Q(
        \input_weight[2][52] ) );
  EDFQD1 \input_weight_reg[2][51]  ( .D(data_in[51]), .E(n491), .CP(clk), .Q(
        \input_weight[2][51] ) );
  EDFQD1 \input_weight_reg[2][50]  ( .D(data_in[50]), .E(n491), .CP(clk), .Q(
        \input_weight[2][50] ) );
  EDFQD1 \input_weight_reg[2][49]  ( .D(data_in[49]), .E(n491), .CP(clk), .Q(
        \input_weight[2][49] ) );
  EDFQD1 \input_weight_reg[2][48]  ( .D(data_in[48]), .E(n491), .CP(clk), .Q(
        \input_weight[2][48] ) );
  EDFQD1 \input_weight_reg[2][47]  ( .D(data_in[47]), .E(n491), .CP(clk), .Q(
        \input_weight[2][47] ) );
  EDFQD1 \input_weight_reg[2][46]  ( .D(data_in[46]), .E(n491), .CP(clk), .Q(
        \input_weight[2][46] ) );
  EDFQD1 \input_weight_reg[2][45]  ( .D(data_in[45]), .E(n491), .CP(clk), .Q(
        \input_weight[2][45] ) );
  EDFQD1 \input_weight_reg[2][44]  ( .D(data_in[44]), .E(n491), .CP(clk), .Q(
        \input_weight[2][44] ) );
  EDFQD1 \input_weight_reg[2][43]  ( .D(data_in[43]), .E(n491), .CP(clk), .Q(
        \input_weight[2][43] ) );
  EDFQD1 \input_weight_reg[2][42]  ( .D(data_in[42]), .E(n491), .CP(clk), .Q(
        \input_weight[2][42] ) );
  EDFQD1 \input_weight_reg[2][41]  ( .D(data_in[41]), .E(n491), .CP(clk), .Q(
        \input_weight[2][41] ) );
  EDFQD1 \input_weight_reg[2][40]  ( .D(data_in[40]), .E(n491), .CP(clk), .Q(
        \input_weight[2][40] ) );
  EDFQD1 \input_weight_reg[2][39]  ( .D(data_in[39]), .E(n491), .CP(clk), .Q(
        \input_weight[2][39] ) );
  EDFQD1 \input_weight_reg[2][38]  ( .D(data_in[38]), .E(n490), .CP(clk), .Q(
        \input_weight[2][38] ) );
  EDFQD1 \input_weight_reg[2][37]  ( .D(data_in[37]), .E(n490), .CP(clk), .Q(
        \input_weight[2][37] ) );
  EDFQD1 \input_weight_reg[2][36]  ( .D(data_in[36]), .E(n490), .CP(clk), .Q(
        \input_weight[2][36] ) );
  EDFQD1 \input_weight_reg[2][35]  ( .D(data_in[35]), .E(n490), .CP(clk), .Q(
        \input_weight[2][35] ) );
  EDFQD1 \input_weight_reg[2][34]  ( .D(data_in[34]), .E(n490), .CP(clk), .Q(
        \input_weight[2][34] ) );
  EDFQD1 \input_weight_reg[2][33]  ( .D(data_in[33]), .E(n490), .CP(clk), .Q(
        \input_weight[2][33] ) );
  EDFQD1 \input_weight_reg[2][32]  ( .D(data_in[32]), .E(n490), .CP(clk), .Q(
        \input_weight[2][32] ) );
  EDFQD1 \input_weight_reg[2][31]  ( .D(data_in[31]), .E(n490), .CP(clk), .Q(
        \input_weight[2][31] ) );
  EDFQD1 \input_weight_reg[2][30]  ( .D(data_in[30]), .E(n490), .CP(clk), .Q(
        \input_weight[2][30] ) );
  EDFQD1 \input_weight_reg[2][29]  ( .D(data_in[29]), .E(n490), .CP(clk), .Q(
        \input_weight[2][29] ) );
  EDFQD1 \input_weight_reg[2][28]  ( .D(data_in[28]), .E(n490), .CP(clk), .Q(
        \input_weight[2][28] ) );
  EDFQD1 \input_weight_reg[2][27]  ( .D(data_in[27]), .E(n490), .CP(clk), .Q(
        \input_weight[2][27] ) );
  EDFQD1 \input_weight_reg[2][26]  ( .D(data_in[26]), .E(n490), .CP(clk), .Q(
        \input_weight[2][26] ) );
  EDFQD1 \input_weight_reg[2][25]  ( .D(data_in[25]), .E(n489), .CP(clk), .Q(
        \input_weight[2][25] ) );
  EDFQD1 \input_weight_reg[2][24]  ( .D(data_in[24]), .E(n489), .CP(clk), .Q(
        \input_weight[2][24] ) );
  EDFQD1 \input_weight_reg[2][23]  ( .D(data_in[23]), .E(n489), .CP(clk), .Q(
        \input_weight[2][23] ) );
  EDFQD1 \input_weight_reg[2][22]  ( .D(data_in[22]), .E(n489), .CP(clk), .Q(
        \input_weight[2][22] ) );
  EDFQD1 \input_weight_reg[2][21]  ( .D(data_in[21]), .E(n489), .CP(clk), .Q(
        \input_weight[2][21] ) );
  EDFQD1 \input_weight_reg[2][20]  ( .D(data_in[20]), .E(n489), .CP(clk), .Q(
        \input_weight[2][20] ) );
  EDFQD1 \input_weight_reg[2][19]  ( .D(data_in[19]), .E(n489), .CP(clk), .Q(
        \input_weight[2][19] ) );
  EDFQD1 \input_weight_reg[2][18]  ( .D(data_in[18]), .E(n489), .CP(clk), .Q(
        \input_weight[2][18] ) );
  EDFQD1 \input_weight_reg[2][17]  ( .D(data_in[17]), .E(n489), .CP(clk), .Q(
        \input_weight[2][17] ) );
  EDFQD1 \input_weight_reg[2][16]  ( .D(data_in[16]), .E(n489), .CP(clk), .Q(
        \input_weight[2][16] ) );
  EDFQD1 \input_weight_reg[2][15]  ( .D(data_in[15]), .E(n489), .CP(clk), .Q(
        \input_weight[2][15] ) );
  EDFQD1 \input_weight_reg[2][14]  ( .D(data_in[14]), .E(n489), .CP(clk), .Q(
        \input_weight[2][14] ) );
  EDFQD1 \input_weight_reg[2][13]  ( .D(data_in[13]), .E(n489), .CP(clk), .Q(
        \input_weight[2][13] ) );
  EDFQD1 \input_weight_reg[2][12]  ( .D(data_in[12]), .E(n488), .CP(clk), .Q(
        \input_weight[2][12] ) );
  EDFQD1 \input_weight_reg[2][11]  ( .D(data_in[11]), .E(n488), .CP(clk), .Q(
        \input_weight[2][11] ) );
  EDFQD1 \input_weight_reg[2][10]  ( .D(data_in[10]), .E(n488), .CP(clk), .Q(
        \input_weight[2][10] ) );
  EDFQD1 \input_weight_reg[2][9]  ( .D(data_in[9]), .E(n488), .CP(clk), .Q(
        \input_weight[2][9] ) );
  EDFQD1 \input_weight_reg[2][8]  ( .D(data_in[8]), .E(n488), .CP(clk), .Q(
        \input_weight[2][8] ) );
  EDFQD1 \input_weight_reg[2][7]  ( .D(data_in[7]), .E(n488), .CP(clk), .Q(
        \input_weight[2][7] ) );
  EDFQD1 \input_weight_reg[2][6]  ( .D(data_in[6]), .E(n488), .CP(clk), .Q(
        \input_weight[2][6] ) );
  EDFQD1 \input_weight_reg[2][5]  ( .D(data_in[5]), .E(n488), .CP(clk), .Q(
        \input_weight[2][5] ) );
  EDFQD1 \input_weight_reg[2][4]  ( .D(data_in[4]), .E(n488), .CP(clk), .Q(
        \input_weight[2][4] ) );
  EDFQD1 \input_weight_reg[2][3]  ( .D(data_in[3]), .E(n488), .CP(clk), .Q(
        \input_weight[2][3] ) );
  EDFQD1 \input_weight_reg[2][2]  ( .D(data_in[2]), .E(n488), .CP(clk), .Q(
        \input_weight[2][2] ) );
  EDFQD1 \input_weight_reg[2][1]  ( .D(data_in[1]), .E(n488), .CP(clk), .Q(
        \input_weight[2][1] ) );
  EDFQD1 \input_weight_reg[2][0]  ( .D(data_in[0]), .E(n488), .CP(clk), .Q(
        \input_weight[2][0] ) );
  EDFQD1 \input_value_reg[0][99]  ( .D(data_in[99]), .E(n407), .CP(clk), .Q(
        \input_value[0][99] ) );
  EDFQD1 \input_value_reg[0][100]  ( .D(data_in[100]), .E(n407), .CP(clk), .Q(
        \input_value[0][100] ) );
  EDFQD1 \input_value_reg[0][101]  ( .D(data_in[101]), .E(n407), .CP(clk), .Q(
        \input_value[0][101] ) );
  EDFQD1 \input_value_reg[0][102]  ( .D(data_in[102]), .E(n407), .CP(clk), .Q(
        \input_value[0][102] ) );
  EDFQD1 \input_value_reg[0][103]  ( .D(data_in[103]), .E(n407), .CP(clk), .Q(
        \input_value[0][103] ) );
  EDFQD1 \input_value_reg[0][104]  ( .D(data_in[104]), .E(n407), .CP(clk), .Q(
        \input_value[0][104] ) );
  EDFQD1 \input_value_reg[0][105]  ( .D(data_in[105]), .E(n407), .CP(clk), .Q(
        \input_value[0][105] ) );
  EDFQD1 \input_value_reg[0][106]  ( .D(data_in[106]), .E(n407), .CP(clk), .Q(
        \input_value[0][106] ) );
  EDFQD1 \input_value_reg[0][107]  ( .D(data_in[107]), .E(n407), .CP(clk), .Q(
        \input_value[0][107] ) );
  EDFQD1 \input_value_reg[0][108]  ( .D(data_in[108]), .E(n407), .CP(clk), .Q(
        \input_value[0][108] ) );
  EDFQD1 \input_value_reg[0][109]  ( .D(data_in[109]), .E(n407), .CP(clk), .Q(
        \input_value[0][109] ) );
  EDFQD1 \input_value_reg[0][110]  ( .D(data_in[110]), .E(n406), .CP(clk), .Q(
        \input_value[0][110] ) );
  EDFQD1 \input_value_reg[0][111]  ( .D(data_in[111]), .E(n406), .CP(clk), .Q(
        \input_value[0][111] ) );
  EDFQD1 \input_value_reg[0][112]  ( .D(data_in[112]), .E(n406), .CP(clk), .Q(
        \input_value[0][112] ) );
  EDFQD1 \input_value_reg[0][113]  ( .D(data_in[113]), .E(n406), .CP(clk), .Q(
        \input_value[0][113] ) );
  EDFQD1 \input_value_reg[0][114]  ( .D(data_in[114]), .E(n406), .CP(clk), .Q(
        \input_value[0][114] ) );
  EDFQD1 \input_value_reg[0][115]  ( .D(data_in[115]), .E(n406), .CP(clk), .Q(
        \input_value[0][115] ) );
  EDFQD1 \input_value_reg[0][116]  ( .D(data_in[116]), .E(n406), .CP(clk), .Q(
        \input_value[0][116] ) );
  EDFQD1 \input_value_reg[0][117]  ( .D(data_in[117]), .E(n406), .CP(clk), .Q(
        \input_value[0][117] ) );
  EDFQD1 \input_value_reg[0][118]  ( .D(data_in[118]), .E(n406), .CP(clk), .Q(
        \input_value[0][118] ) );
  EDFQD1 \input_value_reg[0][119]  ( .D(data_in[119]), .E(n406), .CP(clk), .Q(
        \input_value[0][119] ) );
  EDFQD1 \input_value_reg[0][120]  ( .D(data_in[120]), .E(n406), .CP(clk), .Q(
        \input_value[0][120] ) );
  EDFQD1 \input_value_reg[0][121]  ( .D(data_in[121]), .E(n406), .CP(clk), .Q(
        \input_value[0][121] ) );
  EDFQD1 \input_value_reg[0][122]  ( .D(data_in[122]), .E(n406), .CP(clk), .Q(
        \input_value[0][122] ) );
  EDFQD1 \input_value_reg[0][123]  ( .D(data_in[123]), .E(n405), .CP(clk), .Q(
        \input_value[0][123] ) );
  EDFQD1 \input_value_reg[0][124]  ( .D(data_in[124]), .E(n405), .CP(clk), .Q(
        \input_value[0][124] ) );
  EDFQD1 \input_value_reg[0][125]  ( .D(data_in[125]), .E(n405), .CP(clk), .Q(
        \input_value[0][125] ) );
  EDFQD1 \input_value_reg[0][126]  ( .D(data_in[126]), .E(n405), .CP(clk), .Q(
        \input_value[0][126] ) );
  EDFQD1 \input_value_reg[0][127]  ( .D(data_in[127]), .E(n405), .CP(clk), .Q(
        \input_value[0][127] ) );
  EDFQD1 \input_value_reg[0][98]  ( .D(data_in[98]), .E(n405), .CP(clk), .Q(
        \input_value[0][98] ) );
  EDFQD1 \input_value_reg[0][97]  ( .D(data_in[97]), .E(n405), .CP(clk), .Q(
        \input_value[0][97] ) );
  EDFQD1 \input_value_reg[0][96]  ( .D(data_in[96]), .E(n405), .CP(clk), .Q(
        \input_value[0][96] ) );
  EDFQD1 \input_value_reg[0][95]  ( .D(data_in[95]), .E(n405), .CP(clk), .Q(
        \input_value[0][95] ) );
  EDFQD1 \input_value_reg[0][94]  ( .D(data_in[94]), .E(n405), .CP(clk), .Q(
        \input_value[0][94] ) );
  EDFQD1 \input_value_reg[0][93]  ( .D(data_in[93]), .E(n405), .CP(clk), .Q(
        \input_value[0][93] ) );
  EDFQD1 \input_value_reg[0][92]  ( .D(data_in[92]), .E(n405), .CP(clk), .Q(
        \input_value[0][92] ) );
  EDFQD1 \input_value_reg[0][91]  ( .D(data_in[91]), .E(n405), .CP(clk), .Q(
        \input_value[0][91] ) );
  EDFQD1 \input_value_reg[0][90]  ( .D(data_in[90]), .E(n404), .CP(clk), .Q(
        \input_value[0][90] ) );
  EDFQD1 \input_value_reg[0][89]  ( .D(data_in[89]), .E(n404), .CP(clk), .Q(
        \input_value[0][89] ) );
  EDFQD1 \input_value_reg[0][88]  ( .D(data_in[88]), .E(n404), .CP(clk), .Q(
        \input_value[0][88] ) );
  EDFQD1 \input_value_reg[0][87]  ( .D(data_in[87]), .E(n404), .CP(clk), .Q(
        \input_value[0][87] ) );
  EDFQD1 \input_value_reg[0][86]  ( .D(data_in[86]), .E(n404), .CP(clk), .Q(
        \input_value[0][86] ) );
  EDFQD1 \input_value_reg[0][85]  ( .D(data_in[85]), .E(n404), .CP(clk), .Q(
        \input_value[0][85] ) );
  EDFQD1 \input_value_reg[0][84]  ( .D(data_in[84]), .E(n404), .CP(clk), .Q(
        \input_value[0][84] ) );
  EDFQD1 \input_value_reg[0][83]  ( .D(data_in[83]), .E(n404), .CP(clk), .Q(
        \input_value[0][83] ) );
  EDFQD1 \input_value_reg[0][82]  ( .D(data_in[82]), .E(n404), .CP(clk), .Q(
        \input_value[0][82] ) );
  EDFQD1 \input_value_reg[0][81]  ( .D(data_in[81]), .E(n404), .CP(clk), .Q(
        \input_value[0][81] ) );
  EDFQD1 \input_value_reg[0][80]  ( .D(data_in[80]), .E(n404), .CP(clk), .Q(
        \input_value[0][80] ) );
  EDFQD1 \input_value_reg[0][79]  ( .D(data_in[79]), .E(n404), .CP(clk), .Q(
        \input_value[0][79] ) );
  EDFQD1 \input_value_reg[0][78]  ( .D(data_in[78]), .E(n404), .CP(clk), .Q(
        \input_value[0][78] ) );
  EDFQD1 \input_value_reg[0][77]  ( .D(data_in[77]), .E(n403), .CP(clk), .Q(
        \input_value[0][77] ) );
  EDFQD1 \input_value_reg[0][76]  ( .D(data_in[76]), .E(n403), .CP(clk), .Q(
        \input_value[0][76] ) );
  EDFQD1 \input_value_reg[0][75]  ( .D(data_in[75]), .E(n403), .CP(clk), .Q(
        \input_value[0][75] ) );
  EDFQD1 \input_value_reg[0][74]  ( .D(data_in[74]), .E(n403), .CP(clk), .Q(
        \input_value[0][74] ) );
  EDFQD1 \input_value_reg[0][73]  ( .D(data_in[73]), .E(n403), .CP(clk), .Q(
        \input_value[0][73] ) );
  EDFQD1 \input_value_reg[0][72]  ( .D(data_in[72]), .E(n403), .CP(clk), .Q(
        \input_value[0][72] ) );
  EDFQD1 \input_value_reg[0][71]  ( .D(data_in[71]), .E(n403), .CP(clk), .Q(
        \input_value[0][71] ) );
  EDFQD1 \input_value_reg[0][70]  ( .D(data_in[70]), .E(n403), .CP(clk), .Q(
        \input_value[0][70] ) );
  EDFQD1 \input_value_reg[0][69]  ( .D(data_in[69]), .E(n403), .CP(clk), .Q(
        \input_value[0][69] ) );
  EDFQD1 \input_value_reg[0][68]  ( .D(data_in[68]), .E(n403), .CP(clk), .Q(
        \input_value[0][68] ) );
  EDFQD1 \input_value_reg[0][67]  ( .D(data_in[67]), .E(n403), .CP(clk), .Q(
        \input_value[0][67] ) );
  EDFQD1 \input_value_reg[0][66]  ( .D(data_in[66]), .E(n403), .CP(clk), .Q(
        \input_value[0][66] ) );
  EDFQD1 \input_value_reg[0][65]  ( .D(data_in[65]), .E(n403), .CP(clk), .Q(
        \input_value[0][65] ) );
  EDFQD1 \input_value_reg[0][64]  ( .D(data_in[64]), .E(n402), .CP(clk), .Q(
        \input_value[0][64] ) );
  EDFQD1 \input_value_reg[0][63]  ( .D(data_in[63]), .E(n402), .CP(clk), .Q(
        \input_value[0][63] ) );
  EDFQD1 \input_value_reg[0][62]  ( .D(data_in[62]), .E(n402), .CP(clk), .Q(
        \input_value[0][62] ) );
  EDFQD1 \input_value_reg[0][61]  ( .D(data_in[61]), .E(n402), .CP(clk), .Q(
        \input_value[0][61] ) );
  EDFQD1 \input_value_reg[0][60]  ( .D(data_in[60]), .E(n402), .CP(clk), .Q(
        \input_value[0][60] ) );
  EDFQD1 \input_value_reg[0][59]  ( .D(data_in[59]), .E(n402), .CP(clk), .Q(
        \input_value[0][59] ) );
  EDFQD1 \input_value_reg[0][58]  ( .D(data_in[58]), .E(n402), .CP(clk), .Q(
        \input_value[0][58] ) );
  EDFQD1 \input_value_reg[0][57]  ( .D(data_in[57]), .E(n402), .CP(clk), .Q(
        \input_value[0][57] ) );
  EDFQD1 \input_value_reg[0][56]  ( .D(data_in[56]), .E(n402), .CP(clk), .Q(
        \input_value[0][56] ) );
  EDFQD1 \input_value_reg[0][55]  ( .D(data_in[55]), .E(n402), .CP(clk), .Q(
        \input_value[0][55] ) );
  EDFQD1 \input_value_reg[0][54]  ( .D(data_in[54]), .E(n402), .CP(clk), .Q(
        \input_value[0][54] ) );
  EDFQD1 \input_value_reg[0][53]  ( .D(data_in[53]), .E(n402), .CP(clk), .Q(
        \input_value[0][53] ) );
  EDFQD1 \input_value_reg[0][52]  ( .D(data_in[52]), .E(n402), .CP(clk), .Q(
        \input_value[0][52] ) );
  EDFQD1 \input_value_reg[0][51]  ( .D(data_in[51]), .E(n401), .CP(clk), .Q(
        \input_value[0][51] ) );
  EDFQD1 \input_value_reg[0][50]  ( .D(data_in[50]), .E(n401), .CP(clk), .Q(
        \input_value[0][50] ) );
  EDFQD1 \input_value_reg[0][49]  ( .D(data_in[49]), .E(n401), .CP(clk), .Q(
        \input_value[0][49] ) );
  EDFQD1 \input_value_reg[0][48]  ( .D(data_in[48]), .E(n401), .CP(clk), .Q(
        \input_value[0][48] ) );
  EDFQD1 \input_value_reg[0][47]  ( .D(data_in[47]), .E(n401), .CP(clk), .Q(
        \input_value[0][47] ) );
  EDFQD1 \input_value_reg[0][46]  ( .D(data_in[46]), .E(n401), .CP(clk), .Q(
        \input_value[0][46] ) );
  EDFQD1 \input_value_reg[0][45]  ( .D(data_in[45]), .E(n401), .CP(clk), .Q(
        \input_value[0][45] ) );
  EDFQD1 \input_value_reg[0][44]  ( .D(data_in[44]), .E(n401), .CP(clk), .Q(
        \input_value[0][44] ) );
  EDFQD1 \input_value_reg[0][43]  ( .D(data_in[43]), .E(n401), .CP(clk), .Q(
        \input_value[0][43] ) );
  EDFQD1 \input_value_reg[0][42]  ( .D(data_in[42]), .E(n401), .CP(clk), .Q(
        \input_value[0][42] ) );
  EDFQD1 \input_value_reg[0][41]  ( .D(data_in[41]), .E(n401), .CP(clk), .Q(
        \input_value[0][41] ) );
  EDFQD1 \input_value_reg[0][40]  ( .D(data_in[40]), .E(n401), .CP(clk), .Q(
        \input_value[0][40] ) );
  EDFQD1 \input_value_reg[0][39]  ( .D(data_in[39]), .E(n401), .CP(clk), .Q(
        \input_value[0][39] ) );
  EDFQD1 \input_value_reg[0][38]  ( .D(data_in[38]), .E(n400), .CP(clk), .Q(
        \input_value[0][38] ) );
  EDFQD1 \input_value_reg[0][37]  ( .D(data_in[37]), .E(n400), .CP(clk), .Q(
        \input_value[0][37] ) );
  EDFQD1 \input_value_reg[0][36]  ( .D(data_in[36]), .E(n400), .CP(clk), .Q(
        \input_value[0][36] ) );
  EDFQD1 \input_value_reg[0][35]  ( .D(data_in[35]), .E(n400), .CP(clk), .Q(
        \input_value[0][35] ) );
  EDFQD1 \input_value_reg[0][34]  ( .D(data_in[34]), .E(n400), .CP(clk), .Q(
        \input_value[0][34] ) );
  EDFQD1 \input_value_reg[0][33]  ( .D(data_in[33]), .E(n400), .CP(clk), .Q(
        \input_value[0][33] ) );
  EDFQD1 \input_value_reg[0][32]  ( .D(data_in[32]), .E(n400), .CP(clk), .Q(
        \input_value[0][32] ) );
  EDFQD1 \input_value_reg[0][31]  ( .D(data_in[31]), .E(n400), .CP(clk), .Q(
        \input_value[0][31] ) );
  EDFQD1 \input_value_reg[0][30]  ( .D(data_in[30]), .E(n400), .CP(clk), .Q(
        \input_value[0][30] ) );
  EDFQD1 \input_value_reg[0][29]  ( .D(data_in[29]), .E(n400), .CP(clk), .Q(
        \input_value[0][29] ) );
  EDFQD1 \input_value_reg[0][28]  ( .D(data_in[28]), .E(n400), .CP(clk), .Q(
        \input_value[0][28] ) );
  EDFQD1 \input_value_reg[0][27]  ( .D(data_in[27]), .E(n400), .CP(clk), .Q(
        \input_value[0][27] ) );
  EDFQD1 \input_value_reg[0][26]  ( .D(data_in[26]), .E(n400), .CP(clk), .Q(
        \input_value[0][26] ) );
  EDFQD1 \input_value_reg[0][25]  ( .D(data_in[25]), .E(n399), .CP(clk), .Q(
        \input_value[0][25] ) );
  EDFQD1 \input_value_reg[0][24]  ( .D(data_in[24]), .E(n399), .CP(clk), .Q(
        \input_value[0][24] ) );
  EDFQD1 \input_value_reg[0][23]  ( .D(data_in[23]), .E(n399), .CP(clk), .Q(
        \input_value[0][23] ) );
  EDFQD1 \input_value_reg[0][22]  ( .D(data_in[22]), .E(n399), .CP(clk), .Q(
        \input_value[0][22] ) );
  EDFQD1 \input_value_reg[0][21]  ( .D(data_in[21]), .E(n399), .CP(clk), .Q(
        \input_value[0][21] ) );
  EDFQD1 \input_value_reg[0][20]  ( .D(data_in[20]), .E(n399), .CP(clk), .Q(
        \input_value[0][20] ) );
  EDFQD1 \input_value_reg[0][19]  ( .D(data_in[19]), .E(n399), .CP(clk), .Q(
        \input_value[0][19] ) );
  EDFQD1 \input_value_reg[0][18]  ( .D(data_in[18]), .E(n399), .CP(clk), .Q(
        \input_value[0][18] ) );
  EDFQD1 \input_value_reg[0][17]  ( .D(data_in[17]), .E(n399), .CP(clk), .Q(
        \input_value[0][17] ) );
  EDFQD1 \input_value_reg[0][16]  ( .D(data_in[16]), .E(n399), .CP(clk), .Q(
        \input_value[0][16] ) );
  EDFQD1 \input_value_reg[0][15]  ( .D(data_in[15]), .E(n399), .CP(clk), .Q(
        \input_value[0][15] ) );
  EDFQD1 \input_value_reg[0][14]  ( .D(data_in[14]), .E(n399), .CP(clk), .Q(
        \input_value[0][14] ) );
  EDFQD1 \input_value_reg[0][13]  ( .D(data_in[13]), .E(n399), .CP(clk), .Q(
        \input_value[0][13] ) );
  EDFQD1 \input_value_reg[0][12]  ( .D(data_in[12]), .E(n398), .CP(clk), .Q(
        \input_value[0][12] ) );
  EDFQD1 \input_value_reg[0][11]  ( .D(data_in[11]), .E(n398), .CP(clk), .Q(
        \input_value[0][11] ) );
  EDFQD1 \input_value_reg[0][10]  ( .D(data_in[10]), .E(n398), .CP(clk), .Q(
        \input_value[0][10] ) );
  EDFQD1 \input_value_reg[0][9]  ( .D(data_in[9]), .E(n398), .CP(clk), .Q(
        \input_value[0][9] ) );
  EDFQD1 \input_value_reg[0][8]  ( .D(data_in[8]), .E(n398), .CP(clk), .Q(
        \input_value[0][8] ) );
  EDFQD1 \input_value_reg[0][7]  ( .D(data_in[7]), .E(n398), .CP(clk), .Q(
        \input_value[0][7] ) );
  EDFQD1 \input_value_reg[0][6]  ( .D(data_in[6]), .E(n398), .CP(clk), .Q(
        \input_value[0][6] ) );
  EDFQD1 \input_value_reg[0][5]  ( .D(data_in[5]), .E(n398), .CP(clk), .Q(
        \input_value[0][5] ) );
  EDFQD1 \input_value_reg[0][4]  ( .D(data_in[4]), .E(n398), .CP(clk), .Q(
        \input_value[0][4] ) );
  EDFQD1 \input_value_reg[0][3]  ( .D(data_in[3]), .E(n398), .CP(clk), .Q(
        \input_value[0][3] ) );
  EDFQD1 \input_value_reg[0][2]  ( .D(data_in[2]), .E(n398), .CP(clk), .Q(
        \input_value[0][2] ) );
  EDFQD1 \input_value_reg[0][1]  ( .D(data_in[1]), .E(n398), .CP(clk), .Q(
        \input_value[0][1] ) );
  EDFQD1 \input_value_reg[0][0]  ( .D(data_in[0]), .E(n398), .CP(clk), .Q(
        \input_value[0][0] ) );
  EDFQD1 \input_weight_reg[0][99]  ( .D(data_in[99]), .E(n527), .CP(clk), .Q(
        \input_weight[0][99] ) );
  EDFQD1 \input_weight_reg[0][100]  ( .D(data_in[100]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][100] ) );
  EDFQD1 \input_weight_reg[0][101]  ( .D(data_in[101]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][101] ) );
  EDFQD1 \input_weight_reg[0][102]  ( .D(data_in[102]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][102] ) );
  EDFQD1 \input_weight_reg[0][103]  ( .D(data_in[103]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][103] ) );
  EDFQD1 \input_weight_reg[0][104]  ( .D(data_in[104]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][104] ) );
  EDFQD1 \input_weight_reg[0][105]  ( .D(data_in[105]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][105] ) );
  EDFQD1 \input_weight_reg[0][106]  ( .D(data_in[106]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][106] ) );
  EDFQD1 \input_weight_reg[0][107]  ( .D(data_in[107]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][107] ) );
  EDFQD1 \input_weight_reg[0][108]  ( .D(data_in[108]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][108] ) );
  EDFQD1 \input_weight_reg[0][109]  ( .D(data_in[109]), .E(n527), .CP(clk), 
        .Q(\input_weight[0][109] ) );
  EDFQD1 \input_weight_reg[0][110]  ( .D(data_in[110]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][110] ) );
  EDFQD1 \input_weight_reg[0][111]  ( .D(data_in[111]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][111] ) );
  EDFQD1 \input_weight_reg[0][112]  ( .D(data_in[112]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][112] ) );
  EDFQD1 \input_weight_reg[0][113]  ( .D(data_in[113]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][113] ) );
  EDFQD1 \input_weight_reg[0][114]  ( .D(data_in[114]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][114] ) );
  EDFQD1 \input_weight_reg[0][115]  ( .D(data_in[115]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][115] ) );
  EDFQD1 \input_weight_reg[0][116]  ( .D(data_in[116]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][116] ) );
  EDFQD1 \input_weight_reg[0][117]  ( .D(data_in[117]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][117] ) );
  EDFQD1 \input_weight_reg[0][118]  ( .D(data_in[118]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][118] ) );
  EDFQD1 \input_weight_reg[0][119]  ( .D(data_in[119]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][119] ) );
  EDFQD1 \input_weight_reg[0][120]  ( .D(data_in[120]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][120] ) );
  EDFQD1 \input_weight_reg[0][121]  ( .D(data_in[121]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][121] ) );
  EDFQD1 \input_weight_reg[0][122]  ( .D(data_in[122]), .E(n526), .CP(clk), 
        .Q(\input_weight[0][122] ) );
  EDFQD1 \input_weight_reg[0][123]  ( .D(data_in[123]), .E(n525), .CP(clk), 
        .Q(\input_weight[0][123] ) );
  EDFQD1 \input_weight_reg[0][124]  ( .D(data_in[124]), .E(n525), .CP(clk), 
        .Q(\input_weight[0][124] ) );
  EDFQD1 \input_weight_reg[0][125]  ( .D(data_in[125]), .E(n525), .CP(clk), 
        .Q(\input_weight[0][125] ) );
  EDFQD1 \input_weight_reg[0][126]  ( .D(data_in[126]), .E(n525), .CP(clk), 
        .Q(\input_weight[0][126] ) );
  EDFQD1 \input_weight_reg[0][127]  ( .D(data_in[127]), .E(n525), .CP(clk), 
        .Q(\input_weight[0][127] ) );
  EDFQD1 \input_weight_reg[0][98]  ( .D(data_in[98]), .E(n525), .CP(clk), .Q(
        \input_weight[0][98] ) );
  EDFQD1 \input_weight_reg[0][97]  ( .D(data_in[97]), .E(n525), .CP(clk), .Q(
        \input_weight[0][97] ) );
  EDFQD1 \input_weight_reg[0][96]  ( .D(data_in[96]), .E(n525), .CP(clk), .Q(
        \input_weight[0][96] ) );
  EDFQD1 \input_weight_reg[0][95]  ( .D(data_in[95]), .E(n525), .CP(clk), .Q(
        \input_weight[0][95] ) );
  EDFQD1 \input_weight_reg[0][94]  ( .D(data_in[94]), .E(n525), .CP(clk), .Q(
        \input_weight[0][94] ) );
  EDFQD1 \input_weight_reg[0][93]  ( .D(data_in[93]), .E(n525), .CP(clk), .Q(
        \input_weight[0][93] ) );
  EDFQD1 \input_weight_reg[0][92]  ( .D(data_in[92]), .E(n525), .CP(clk), .Q(
        \input_weight[0][92] ) );
  EDFQD1 \input_weight_reg[0][91]  ( .D(data_in[91]), .E(n525), .CP(clk), .Q(
        \input_weight[0][91] ) );
  EDFQD1 \input_weight_reg[0][90]  ( .D(data_in[90]), .E(n524), .CP(clk), .Q(
        \input_weight[0][90] ) );
  EDFQD1 \input_weight_reg[0][89]  ( .D(data_in[89]), .E(n524), .CP(clk), .Q(
        \input_weight[0][89] ) );
  EDFQD1 \input_weight_reg[0][88]  ( .D(data_in[88]), .E(n524), .CP(clk), .Q(
        \input_weight[0][88] ) );
  EDFQD1 \input_weight_reg[0][87]  ( .D(data_in[87]), .E(n524), .CP(clk), .Q(
        \input_weight[0][87] ) );
  EDFQD1 \input_weight_reg[0][86]  ( .D(data_in[86]), .E(n524), .CP(clk), .Q(
        \input_weight[0][86] ) );
  EDFQD1 \input_weight_reg[0][85]  ( .D(data_in[85]), .E(n524), .CP(clk), .Q(
        \input_weight[0][85] ) );
  EDFQD1 \input_weight_reg[0][84]  ( .D(data_in[84]), .E(n524), .CP(clk), .Q(
        \input_weight[0][84] ) );
  EDFQD1 \input_weight_reg[0][83]  ( .D(data_in[83]), .E(n524), .CP(clk), .Q(
        \input_weight[0][83] ) );
  EDFQD1 \input_weight_reg[0][82]  ( .D(data_in[82]), .E(n524), .CP(clk), .Q(
        \input_weight[0][82] ) );
  EDFQD1 \input_weight_reg[0][81]  ( .D(data_in[81]), .E(n524), .CP(clk), .Q(
        \input_weight[0][81] ) );
  EDFQD1 \input_weight_reg[0][80]  ( .D(data_in[80]), .E(n524), .CP(clk), .Q(
        \input_weight[0][80] ) );
  EDFQD1 \input_weight_reg[0][79]  ( .D(data_in[79]), .E(n524), .CP(clk), .Q(
        \input_weight[0][79] ) );
  EDFQD1 \input_weight_reg[0][78]  ( .D(data_in[78]), .E(n524), .CP(clk), .Q(
        \input_weight[0][78] ) );
  EDFQD1 \input_weight_reg[0][77]  ( .D(data_in[77]), .E(n523), .CP(clk), .Q(
        \input_weight[0][77] ) );
  EDFQD1 \input_weight_reg[0][76]  ( .D(data_in[76]), .E(n523), .CP(clk), .Q(
        \input_weight[0][76] ) );
  EDFQD1 \input_weight_reg[0][75]  ( .D(data_in[75]), .E(n523), .CP(clk), .Q(
        \input_weight[0][75] ) );
  EDFQD1 \input_weight_reg[0][74]  ( .D(data_in[74]), .E(n523), .CP(clk), .Q(
        \input_weight[0][74] ) );
  EDFQD1 \input_weight_reg[0][73]  ( .D(data_in[73]), .E(n523), .CP(clk), .Q(
        \input_weight[0][73] ) );
  EDFQD1 \input_weight_reg[0][72]  ( .D(data_in[72]), .E(n523), .CP(clk), .Q(
        \input_weight[0][72] ) );
  EDFQD1 \input_weight_reg[0][71]  ( .D(data_in[71]), .E(n523), .CP(clk), .Q(
        \input_weight[0][71] ) );
  EDFQD1 \input_weight_reg[0][70]  ( .D(data_in[70]), .E(n523), .CP(clk), .Q(
        \input_weight[0][70] ) );
  EDFQD1 \input_weight_reg[0][69]  ( .D(data_in[69]), .E(n523), .CP(clk), .Q(
        \input_weight[0][69] ) );
  EDFQD1 \input_weight_reg[0][68]  ( .D(data_in[68]), .E(n523), .CP(clk), .Q(
        \input_weight[0][68] ) );
  EDFQD1 \input_weight_reg[0][67]  ( .D(data_in[67]), .E(n523), .CP(clk), .Q(
        \input_weight[0][67] ) );
  EDFQD1 \input_weight_reg[0][66]  ( .D(data_in[66]), .E(n523), .CP(clk), .Q(
        \input_weight[0][66] ) );
  EDFQD1 \input_weight_reg[0][65]  ( .D(data_in[65]), .E(n523), .CP(clk), .Q(
        \input_weight[0][65] ) );
  EDFQD1 \input_weight_reg[0][64]  ( .D(data_in[64]), .E(n522), .CP(clk), .Q(
        \input_weight[0][64] ) );
  EDFQD1 \input_weight_reg[0][63]  ( .D(data_in[63]), .E(n522), .CP(clk), .Q(
        \input_weight[0][63] ) );
  EDFQD1 \input_weight_reg[0][62]  ( .D(data_in[62]), .E(n522), .CP(clk), .Q(
        \input_weight[0][62] ) );
  EDFQD1 \input_weight_reg[0][61]  ( .D(data_in[61]), .E(n522), .CP(clk), .Q(
        \input_weight[0][61] ) );
  EDFQD1 \input_weight_reg[0][60]  ( .D(data_in[60]), .E(n522), .CP(clk), .Q(
        \input_weight[0][60] ) );
  EDFQD1 \input_weight_reg[0][59]  ( .D(data_in[59]), .E(n522), .CP(clk), .Q(
        \input_weight[0][59] ) );
  EDFQD1 \input_weight_reg[0][58]  ( .D(data_in[58]), .E(n522), .CP(clk), .Q(
        \input_weight[0][58] ) );
  EDFQD1 \input_weight_reg[0][57]  ( .D(data_in[57]), .E(n522), .CP(clk), .Q(
        \input_weight[0][57] ) );
  EDFQD1 \input_weight_reg[0][56]  ( .D(data_in[56]), .E(n522), .CP(clk), .Q(
        \input_weight[0][56] ) );
  EDFQD1 \input_weight_reg[0][55]  ( .D(data_in[55]), .E(n522), .CP(clk), .Q(
        \input_weight[0][55] ) );
  EDFQD1 \input_weight_reg[0][54]  ( .D(data_in[54]), .E(n522), .CP(clk), .Q(
        \input_weight[0][54] ) );
  EDFQD1 \input_weight_reg[0][53]  ( .D(data_in[53]), .E(n522), .CP(clk), .Q(
        \input_weight[0][53] ) );
  EDFQD1 \input_weight_reg[0][52]  ( .D(data_in[52]), .E(n522), .CP(clk), .Q(
        \input_weight[0][52] ) );
  EDFQD1 \input_weight_reg[0][51]  ( .D(data_in[51]), .E(n521), .CP(clk), .Q(
        \input_weight[0][51] ) );
  EDFQD1 \input_weight_reg[0][50]  ( .D(data_in[50]), .E(n521), .CP(clk), .Q(
        \input_weight[0][50] ) );
  EDFQD1 \input_weight_reg[0][49]  ( .D(data_in[49]), .E(n521), .CP(clk), .Q(
        \input_weight[0][49] ) );
  EDFQD1 \input_weight_reg[0][48]  ( .D(data_in[48]), .E(n521), .CP(clk), .Q(
        \input_weight[0][48] ) );
  EDFQD1 \input_weight_reg[0][47]  ( .D(data_in[47]), .E(n521), .CP(clk), .Q(
        \input_weight[0][47] ) );
  EDFQD1 \input_weight_reg[0][46]  ( .D(data_in[46]), .E(n521), .CP(clk), .Q(
        \input_weight[0][46] ) );
  EDFQD1 \input_weight_reg[0][45]  ( .D(data_in[45]), .E(n521), .CP(clk), .Q(
        \input_weight[0][45] ) );
  EDFQD1 \input_weight_reg[0][44]  ( .D(data_in[44]), .E(n521), .CP(clk), .Q(
        \input_weight[0][44] ) );
  EDFQD1 \input_weight_reg[0][43]  ( .D(data_in[43]), .E(n521), .CP(clk), .Q(
        \input_weight[0][43] ) );
  EDFQD1 \input_weight_reg[0][42]  ( .D(data_in[42]), .E(n521), .CP(clk), .Q(
        \input_weight[0][42] ) );
  EDFQD1 \input_weight_reg[0][41]  ( .D(data_in[41]), .E(n521), .CP(clk), .Q(
        \input_weight[0][41] ) );
  EDFQD1 \input_weight_reg[0][40]  ( .D(data_in[40]), .E(n521), .CP(clk), .Q(
        \input_weight[0][40] ) );
  EDFQD1 \input_weight_reg[0][39]  ( .D(data_in[39]), .E(n521), .CP(clk), .Q(
        \input_weight[0][39] ) );
  EDFQD1 \input_weight_reg[0][38]  ( .D(data_in[38]), .E(n520), .CP(clk), .Q(
        \input_weight[0][38] ) );
  EDFQD1 \input_weight_reg[0][37]  ( .D(data_in[37]), .E(n520), .CP(clk), .Q(
        \input_weight[0][37] ) );
  EDFQD1 \input_weight_reg[0][36]  ( .D(data_in[36]), .E(n520), .CP(clk), .Q(
        \input_weight[0][36] ) );
  EDFQD1 \input_weight_reg[0][35]  ( .D(data_in[35]), .E(n520), .CP(clk), .Q(
        \input_weight[0][35] ) );
  EDFQD1 \input_weight_reg[0][34]  ( .D(data_in[34]), .E(n520), .CP(clk), .Q(
        \input_weight[0][34] ) );
  EDFQD1 \input_weight_reg[0][33]  ( .D(data_in[33]), .E(n520), .CP(clk), .Q(
        \input_weight[0][33] ) );
  EDFQD1 \input_weight_reg[0][32]  ( .D(data_in[32]), .E(n520), .CP(clk), .Q(
        \input_weight[0][32] ) );
  EDFQD1 \input_weight_reg[0][31]  ( .D(data_in[31]), .E(n520), .CP(clk), .Q(
        \input_weight[0][31] ) );
  EDFQD1 \input_weight_reg[0][30]  ( .D(data_in[30]), .E(n520), .CP(clk), .Q(
        \input_weight[0][30] ) );
  EDFQD1 \input_weight_reg[0][29]  ( .D(data_in[29]), .E(n520), .CP(clk), .Q(
        \input_weight[0][29] ) );
  EDFQD1 \input_weight_reg[0][28]  ( .D(data_in[28]), .E(n520), .CP(clk), .Q(
        \input_weight[0][28] ) );
  EDFQD1 \input_weight_reg[0][27]  ( .D(data_in[27]), .E(n520), .CP(clk), .Q(
        \input_weight[0][27] ) );
  EDFQD1 \input_weight_reg[0][26]  ( .D(data_in[26]), .E(n520), .CP(clk), .Q(
        \input_weight[0][26] ) );
  EDFQD1 \input_weight_reg[0][25]  ( .D(data_in[25]), .E(n519), .CP(clk), .Q(
        \input_weight[0][25] ) );
  EDFQD1 \input_weight_reg[0][24]  ( .D(data_in[24]), .E(n519), .CP(clk), .Q(
        \input_weight[0][24] ) );
  EDFQD1 \input_weight_reg[0][23]  ( .D(data_in[23]), .E(n519), .CP(clk), .Q(
        \input_weight[0][23] ) );
  EDFQD1 \input_weight_reg[0][22]  ( .D(data_in[22]), .E(n519), .CP(clk), .Q(
        \input_weight[0][22] ) );
  EDFQD1 \input_weight_reg[0][21]  ( .D(data_in[21]), .E(n519), .CP(clk), .Q(
        \input_weight[0][21] ) );
  EDFQD1 \input_weight_reg[0][20]  ( .D(data_in[20]), .E(n519), .CP(clk), .Q(
        \input_weight[0][20] ) );
  EDFQD1 \input_weight_reg[0][19]  ( .D(data_in[19]), .E(n519), .CP(clk), .Q(
        \input_weight[0][19] ) );
  EDFQD1 \input_weight_reg[0][18]  ( .D(data_in[18]), .E(n519), .CP(clk), .Q(
        \input_weight[0][18] ) );
  EDFQD1 \input_weight_reg[0][17]  ( .D(data_in[17]), .E(n519), .CP(clk), .Q(
        \input_weight[0][17] ) );
  EDFQD1 \input_weight_reg[0][16]  ( .D(data_in[16]), .E(n519), .CP(clk), .Q(
        \input_weight[0][16] ) );
  EDFQD1 \input_weight_reg[0][15]  ( .D(data_in[15]), .E(n519), .CP(clk), .Q(
        \input_weight[0][15] ) );
  EDFQD1 \input_weight_reg[0][14]  ( .D(data_in[14]), .E(n519), .CP(clk), .Q(
        \input_weight[0][14] ) );
  EDFQD1 \input_weight_reg[0][13]  ( .D(data_in[13]), .E(n519), .CP(clk), .Q(
        \input_weight[0][13] ) );
  EDFQD1 \input_weight_reg[0][12]  ( .D(data_in[12]), .E(n518), .CP(clk), .Q(
        \input_weight[0][12] ) );
  EDFQD1 \input_weight_reg[0][11]  ( .D(data_in[11]), .E(n518), .CP(clk), .Q(
        \input_weight[0][11] ) );
  EDFQD1 \input_weight_reg[0][10]  ( .D(data_in[10]), .E(n518), .CP(clk), .Q(
        \input_weight[0][10] ) );
  EDFQD1 \input_weight_reg[0][9]  ( .D(data_in[9]), .E(n518), .CP(clk), .Q(
        \input_weight[0][9] ) );
  EDFQD1 \input_weight_reg[0][8]  ( .D(data_in[8]), .E(n518), .CP(clk), .Q(
        \input_weight[0][8] ) );
  EDFQD1 \input_weight_reg[0][7]  ( .D(data_in[7]), .E(n518), .CP(clk), .Q(
        \input_weight[0][7] ) );
  EDFQD1 \input_weight_reg[0][6]  ( .D(data_in[6]), .E(n518), .CP(clk), .Q(
        \input_weight[0][6] ) );
  EDFQD1 \input_weight_reg[0][5]  ( .D(data_in[5]), .E(n518), .CP(clk), .Q(
        \input_weight[0][5] ) );
  EDFQD1 \input_weight_reg[0][4]  ( .D(data_in[4]), .E(n518), .CP(clk), .Q(
        \input_weight[0][4] ) );
  EDFQD1 \input_weight_reg[0][3]  ( .D(data_in[3]), .E(n518), .CP(clk), .Q(
        \input_weight[0][3] ) );
  EDFQD1 \input_weight_reg[0][2]  ( .D(data_in[2]), .E(n518), .CP(clk), .Q(
        \input_weight[0][2] ) );
  EDFQD1 \input_weight_reg[0][1]  ( .D(data_in[1]), .E(n518), .CP(clk), .Q(
        \input_weight[0][1] ) );
  EDFQD1 \input_weight_reg[0][0]  ( .D(data_in[0]), .E(n518), .CP(clk), .Q(
        \input_weight[0][0] ) );
  EDFQD1 \input_value_reg[7][99]  ( .D(data_in[99]), .E(n302), .CP(clk), .Q(
        \input_value[7][99] ) );
  EDFQD1 \input_value_reg[7][100]  ( .D(data_in[100]), .E(n302), .CP(clk), .Q(
        \input_value[7][100] ) );
  EDFQD1 \input_value_reg[7][101]  ( .D(data_in[101]), .E(n302), .CP(clk), .Q(
        \input_value[7][101] ) );
  EDFQD1 \input_value_reg[7][102]  ( .D(data_in[102]), .E(n302), .CP(clk), .Q(
        \input_value[7][102] ) );
  EDFQD1 \input_value_reg[7][103]  ( .D(data_in[103]), .E(n302), .CP(clk), .Q(
        \input_value[7][103] ) );
  EDFQD1 \input_value_reg[7][104]  ( .D(data_in[104]), .E(n302), .CP(clk), .Q(
        \input_value[7][104] ) );
  EDFQD1 \input_value_reg[7][105]  ( .D(data_in[105]), .E(n302), .CP(clk), .Q(
        \input_value[7][105] ) );
  EDFQD1 \input_value_reg[7][106]  ( .D(data_in[106]), .E(n302), .CP(clk), .Q(
        \input_value[7][106] ) );
  EDFQD1 \input_value_reg[7][107]  ( .D(data_in[107]), .E(n302), .CP(clk), .Q(
        \input_value[7][107] ) );
  EDFQD1 \input_value_reg[7][108]  ( .D(data_in[108]), .E(n302), .CP(clk), .Q(
        \input_value[7][108] ) );
  EDFQD1 \input_value_reg[7][109]  ( .D(data_in[109]), .E(n302), .CP(clk), .Q(
        \input_value[7][109] ) );
  EDFQD1 \input_value_reg[7][110]  ( .D(data_in[110]), .E(n301), .CP(clk), .Q(
        \input_value[7][110] ) );
  EDFQD1 \input_value_reg[7][111]  ( .D(data_in[111]), .E(n301), .CP(clk), .Q(
        \input_value[7][111] ) );
  EDFQD1 \input_value_reg[7][112]  ( .D(data_in[112]), .E(n301), .CP(clk), .Q(
        \input_value[7][112] ) );
  EDFQD1 \input_value_reg[7][113]  ( .D(data_in[113]), .E(n301), .CP(clk), .Q(
        \input_value[7][113] ) );
  EDFQD1 \input_value_reg[7][114]  ( .D(data_in[114]), .E(n301), .CP(clk), .Q(
        \input_value[7][114] ) );
  EDFQD1 \input_value_reg[7][115]  ( .D(data_in[115]), .E(n301), .CP(clk), .Q(
        \input_value[7][115] ) );
  EDFQD1 \input_value_reg[7][116]  ( .D(data_in[116]), .E(n301), .CP(clk), .Q(
        \input_value[7][116] ) );
  EDFQD1 \input_value_reg[7][117]  ( .D(data_in[117]), .E(n301), .CP(clk), .Q(
        \input_value[7][117] ) );
  EDFQD1 \input_value_reg[7][118]  ( .D(data_in[118]), .E(n301), .CP(clk), .Q(
        \input_value[7][118] ) );
  EDFQD1 \input_value_reg[7][119]  ( .D(data_in[119]), .E(n301), .CP(clk), .Q(
        \input_value[7][119] ) );
  EDFQD1 \input_value_reg[7][120]  ( .D(data_in[120]), .E(n301), .CP(clk), .Q(
        \input_value[7][120] ) );
  EDFQD1 \input_value_reg[7][121]  ( .D(data_in[121]), .E(n301), .CP(clk), .Q(
        \input_value[7][121] ) );
  EDFQD1 \input_value_reg[7][122]  ( .D(data_in[122]), .E(n301), .CP(clk), .Q(
        \input_value[7][122] ) );
  EDFQD1 \input_value_reg[7][123]  ( .D(data_in[123]), .E(n300), .CP(clk), .Q(
        \input_value[7][123] ) );
  EDFQD1 \input_value_reg[7][124]  ( .D(data_in[124]), .E(n300), .CP(clk), .Q(
        \input_value[7][124] ) );
  EDFQD1 \input_value_reg[7][125]  ( .D(data_in[125]), .E(n300), .CP(clk), .Q(
        \input_value[7][125] ) );
  EDFQD1 \input_value_reg[7][126]  ( .D(data_in[126]), .E(n300), .CP(clk), .Q(
        \input_value[7][126] ) );
  EDFQD1 \input_value_reg[7][127]  ( .D(data_in[127]), .E(n300), .CP(clk), .Q(
        \input_value[7][127] ) );
  EDFQD1 \input_value_reg[7][98]  ( .D(data_in[98]), .E(n300), .CP(clk), .Q(
        \input_value[7][98] ) );
  EDFQD1 \input_value_reg[7][97]  ( .D(data_in[97]), .E(n300), .CP(clk), .Q(
        \input_value[7][97] ) );
  EDFQD1 \input_value_reg[7][96]  ( .D(data_in[96]), .E(n300), .CP(clk), .Q(
        \input_value[7][96] ) );
  EDFQD1 \input_value_reg[7][95]  ( .D(data_in[95]), .E(n300), .CP(clk), .Q(
        \input_value[7][95] ) );
  EDFQD1 \input_value_reg[7][94]  ( .D(data_in[94]), .E(n300), .CP(clk), .Q(
        \input_value[7][94] ) );
  EDFQD1 \input_value_reg[7][93]  ( .D(data_in[93]), .E(n300), .CP(clk), .Q(
        \input_value[7][93] ) );
  EDFQD1 \input_value_reg[7][92]  ( .D(data_in[92]), .E(n300), .CP(clk), .Q(
        \input_value[7][92] ) );
  EDFQD1 \input_value_reg[7][91]  ( .D(data_in[91]), .E(n300), .CP(clk), .Q(
        \input_value[7][91] ) );
  EDFQD1 \input_value_reg[7][90]  ( .D(data_in[90]), .E(n299), .CP(clk), .Q(
        \input_value[7][90] ) );
  EDFQD1 \input_value_reg[7][89]  ( .D(data_in[89]), .E(n299), .CP(clk), .Q(
        \input_value[7][89] ) );
  EDFQD1 \input_value_reg[7][88]  ( .D(data_in[88]), .E(n299), .CP(clk), .Q(
        \input_value[7][88] ) );
  EDFQD1 \input_value_reg[7][87]  ( .D(data_in[87]), .E(n299), .CP(clk), .Q(
        \input_value[7][87] ) );
  EDFQD1 \input_value_reg[7][86]  ( .D(data_in[86]), .E(n299), .CP(clk), .Q(
        \input_value[7][86] ) );
  EDFQD1 \input_value_reg[7][85]  ( .D(data_in[85]), .E(n299), .CP(clk), .Q(
        \input_value[7][85] ) );
  EDFQD1 \input_value_reg[7][84]  ( .D(data_in[84]), .E(n299), .CP(clk), .Q(
        \input_value[7][84] ) );
  EDFQD1 \input_value_reg[7][83]  ( .D(data_in[83]), .E(n299), .CP(clk), .Q(
        \input_value[7][83] ) );
  EDFQD1 \input_value_reg[7][82]  ( .D(data_in[82]), .E(n299), .CP(clk), .Q(
        \input_value[7][82] ) );
  EDFQD1 \input_value_reg[7][81]  ( .D(data_in[81]), .E(n299), .CP(clk), .Q(
        \input_value[7][81] ) );
  EDFQD1 \input_value_reg[7][80]  ( .D(data_in[80]), .E(n299), .CP(clk), .Q(
        \input_value[7][80] ) );
  EDFQD1 \input_value_reg[7][79]  ( .D(data_in[79]), .E(n299), .CP(clk), .Q(
        \input_value[7][79] ) );
  EDFQD1 \input_value_reg[7][78]  ( .D(data_in[78]), .E(n299), .CP(clk), .Q(
        \input_value[7][78] ) );
  EDFQD1 \input_value_reg[7][77]  ( .D(data_in[77]), .E(n298), .CP(clk), .Q(
        \input_value[7][77] ) );
  EDFQD1 \input_value_reg[7][76]  ( .D(data_in[76]), .E(n298), .CP(clk), .Q(
        \input_value[7][76] ) );
  EDFQD1 \input_value_reg[7][75]  ( .D(data_in[75]), .E(n298), .CP(clk), .Q(
        \input_value[7][75] ) );
  EDFQD1 \input_value_reg[7][74]  ( .D(data_in[74]), .E(n298), .CP(clk), .Q(
        \input_value[7][74] ) );
  EDFQD1 \input_value_reg[7][73]  ( .D(data_in[73]), .E(n298), .CP(clk), .Q(
        \input_value[7][73] ) );
  EDFQD1 \input_value_reg[7][72]  ( .D(data_in[72]), .E(n298), .CP(clk), .Q(
        \input_value[7][72] ) );
  EDFQD1 \input_value_reg[7][71]  ( .D(data_in[71]), .E(n298), .CP(clk), .Q(
        \input_value[7][71] ) );
  EDFQD1 \input_value_reg[7][70]  ( .D(data_in[70]), .E(n298), .CP(clk), .Q(
        \input_value[7][70] ) );
  EDFQD1 \input_value_reg[7][69]  ( .D(data_in[69]), .E(n298), .CP(clk), .Q(
        \input_value[7][69] ) );
  EDFQD1 \input_value_reg[7][68]  ( .D(data_in[68]), .E(n298), .CP(clk), .Q(
        \input_value[7][68] ) );
  EDFQD1 \input_value_reg[7][67]  ( .D(data_in[67]), .E(n298), .CP(clk), .Q(
        \input_value[7][67] ) );
  EDFQD1 \input_value_reg[7][66]  ( .D(data_in[66]), .E(n298), .CP(clk), .Q(
        \input_value[7][66] ) );
  EDFQD1 \input_value_reg[7][65]  ( .D(data_in[65]), .E(n298), .CP(clk), .Q(
        \input_value[7][65] ) );
  EDFQD1 \input_value_reg[7][64]  ( .D(data_in[64]), .E(n297), .CP(clk), .Q(
        \input_value[7][64] ) );
  EDFQD1 \input_value_reg[7][63]  ( .D(data_in[63]), .E(n297), .CP(clk), .Q(
        \input_value[7][63] ) );
  EDFQD1 \input_value_reg[7][62]  ( .D(data_in[62]), .E(n297), .CP(clk), .Q(
        \input_value[7][62] ) );
  EDFQD1 \input_value_reg[7][61]  ( .D(data_in[61]), .E(n297), .CP(clk), .Q(
        \input_value[7][61] ) );
  EDFQD1 \input_value_reg[7][60]  ( .D(data_in[60]), .E(n297), .CP(clk), .Q(
        \input_value[7][60] ) );
  EDFQD1 \input_value_reg[7][59]  ( .D(data_in[59]), .E(n297), .CP(clk), .Q(
        \input_value[7][59] ) );
  EDFQD1 \input_value_reg[7][58]  ( .D(data_in[58]), .E(n297), .CP(clk), .Q(
        \input_value[7][58] ) );
  EDFQD1 \input_value_reg[7][57]  ( .D(data_in[57]), .E(n297), .CP(clk), .Q(
        \input_value[7][57] ) );
  EDFQD1 \input_value_reg[7][56]  ( .D(data_in[56]), .E(n297), .CP(clk), .Q(
        \input_value[7][56] ) );
  EDFQD1 \input_value_reg[7][55]  ( .D(data_in[55]), .E(n297), .CP(clk), .Q(
        \input_value[7][55] ) );
  EDFQD1 \input_value_reg[7][54]  ( .D(data_in[54]), .E(n297), .CP(clk), .Q(
        \input_value[7][54] ) );
  EDFQD1 \input_value_reg[7][53]  ( .D(data_in[53]), .E(n297), .CP(clk), .Q(
        \input_value[7][53] ) );
  EDFQD1 \input_value_reg[7][52]  ( .D(data_in[52]), .E(n297), .CP(clk), .Q(
        \input_value[7][52] ) );
  EDFQD1 \input_value_reg[7][51]  ( .D(data_in[51]), .E(n296), .CP(clk), .Q(
        \input_value[7][51] ) );
  EDFQD1 \input_value_reg[7][50]  ( .D(data_in[50]), .E(n296), .CP(clk), .Q(
        \input_value[7][50] ) );
  EDFQD1 \input_value_reg[7][49]  ( .D(data_in[49]), .E(n296), .CP(clk), .Q(
        \input_value[7][49] ) );
  EDFQD1 \input_value_reg[7][48]  ( .D(data_in[48]), .E(n296), .CP(clk), .Q(
        \input_value[7][48] ) );
  EDFQD1 \input_value_reg[7][47]  ( .D(data_in[47]), .E(n296), .CP(clk), .Q(
        \input_value[7][47] ) );
  EDFQD1 \input_value_reg[7][46]  ( .D(data_in[46]), .E(n296), .CP(clk), .Q(
        \input_value[7][46] ) );
  EDFQD1 \input_value_reg[7][45]  ( .D(data_in[45]), .E(n296), .CP(clk), .Q(
        \input_value[7][45] ) );
  EDFQD1 \input_value_reg[7][44]  ( .D(data_in[44]), .E(n296), .CP(clk), .Q(
        \input_value[7][44] ) );
  EDFQD1 \input_value_reg[7][43]  ( .D(data_in[43]), .E(n296), .CP(clk), .Q(
        \input_value[7][43] ) );
  EDFQD1 \input_value_reg[7][42]  ( .D(data_in[42]), .E(n296), .CP(clk), .Q(
        \input_value[7][42] ) );
  EDFQD1 \input_value_reg[7][41]  ( .D(data_in[41]), .E(n296), .CP(clk), .Q(
        \input_value[7][41] ) );
  EDFQD1 \input_value_reg[7][40]  ( .D(data_in[40]), .E(n296), .CP(clk), .Q(
        \input_value[7][40] ) );
  EDFQD1 \input_value_reg[7][39]  ( .D(data_in[39]), .E(n296), .CP(clk), .Q(
        \input_value[7][39] ) );
  EDFQD1 \input_value_reg[7][38]  ( .D(data_in[38]), .E(n295), .CP(clk), .Q(
        \input_value[7][38] ) );
  EDFQD1 \input_value_reg[7][37]  ( .D(data_in[37]), .E(n295), .CP(clk), .Q(
        \input_value[7][37] ) );
  EDFQD1 \input_value_reg[7][36]  ( .D(data_in[36]), .E(n295), .CP(clk), .Q(
        \input_value[7][36] ) );
  EDFQD1 \input_value_reg[7][35]  ( .D(data_in[35]), .E(n295), .CP(clk), .Q(
        \input_value[7][35] ) );
  EDFQD1 \input_value_reg[7][34]  ( .D(data_in[34]), .E(n295), .CP(clk), .Q(
        \input_value[7][34] ) );
  EDFQD1 \input_value_reg[7][33]  ( .D(data_in[33]), .E(n295), .CP(clk), .Q(
        \input_value[7][33] ) );
  EDFQD1 \input_value_reg[7][32]  ( .D(data_in[32]), .E(n295), .CP(clk), .Q(
        \input_value[7][32] ) );
  EDFQD1 \input_value_reg[7][31]  ( .D(data_in[31]), .E(n295), .CP(clk), .Q(
        \input_value[7][31] ) );
  EDFQD1 \input_value_reg[7][30]  ( .D(data_in[30]), .E(n295), .CP(clk), .Q(
        \input_value[7][30] ) );
  EDFQD1 \input_value_reg[7][29]  ( .D(data_in[29]), .E(n295), .CP(clk), .Q(
        \input_value[7][29] ) );
  EDFQD1 \input_value_reg[7][28]  ( .D(data_in[28]), .E(n295), .CP(clk), .Q(
        \input_value[7][28] ) );
  EDFQD1 \input_value_reg[7][27]  ( .D(data_in[27]), .E(n295), .CP(clk), .Q(
        \input_value[7][27] ) );
  EDFQD1 \input_value_reg[7][26]  ( .D(data_in[26]), .E(n295), .CP(clk), .Q(
        \input_value[7][26] ) );
  EDFQD1 \input_value_reg[7][25]  ( .D(data_in[25]), .E(n294), .CP(clk), .Q(
        \input_value[7][25] ) );
  EDFQD1 \input_value_reg[7][24]  ( .D(data_in[24]), .E(n294), .CP(clk), .Q(
        \input_value[7][24] ) );
  EDFQD1 \input_value_reg[7][23]  ( .D(data_in[23]), .E(n294), .CP(clk), .Q(
        \input_value[7][23] ) );
  EDFQD1 \input_value_reg[7][22]  ( .D(data_in[22]), .E(n294), .CP(clk), .Q(
        \input_value[7][22] ) );
  EDFQD1 \input_value_reg[7][21]  ( .D(data_in[21]), .E(n294), .CP(clk), .Q(
        \input_value[7][21] ) );
  EDFQD1 \input_value_reg[7][20]  ( .D(data_in[20]), .E(n294), .CP(clk), .Q(
        \input_value[7][20] ) );
  EDFQD1 \input_value_reg[7][19]  ( .D(data_in[19]), .E(n294), .CP(clk), .Q(
        \input_value[7][19] ) );
  EDFQD1 \input_value_reg[7][18]  ( .D(data_in[18]), .E(n294), .CP(clk), .Q(
        \input_value[7][18] ) );
  EDFQD1 \input_value_reg[7][17]  ( .D(data_in[17]), .E(n294), .CP(clk), .Q(
        \input_value[7][17] ) );
  EDFQD1 \input_value_reg[7][16]  ( .D(data_in[16]), .E(n294), .CP(clk), .Q(
        \input_value[7][16] ) );
  EDFQD1 \input_value_reg[7][15]  ( .D(data_in[15]), .E(n294), .CP(clk), .Q(
        \input_value[7][15] ) );
  EDFQD1 \input_value_reg[7][14]  ( .D(data_in[14]), .E(n294), .CP(clk), .Q(
        \input_value[7][14] ) );
  EDFQD1 \input_value_reg[7][13]  ( .D(data_in[13]), .E(n294), .CP(clk), .Q(
        \input_value[7][13] ) );
  EDFQD1 \input_value_reg[7][12]  ( .D(data_in[12]), .E(n293), .CP(clk), .Q(
        \input_value[7][12] ) );
  EDFQD1 \input_value_reg[7][11]  ( .D(data_in[11]), .E(n293), .CP(clk), .Q(
        \input_value[7][11] ) );
  EDFQD1 \input_value_reg[7][10]  ( .D(data_in[10]), .E(n293), .CP(clk), .Q(
        \input_value[7][10] ) );
  EDFQD1 \input_value_reg[7][9]  ( .D(data_in[9]), .E(n293), .CP(clk), .Q(
        \input_value[7][9] ) );
  EDFQD1 \input_value_reg[7][8]  ( .D(data_in[8]), .E(n293), .CP(clk), .Q(
        \input_value[7][8] ) );
  EDFQD1 \input_value_reg[7][7]  ( .D(data_in[7]), .E(n293), .CP(clk), .Q(
        \input_value[7][7] ) );
  EDFQD1 \input_value_reg[7][6]  ( .D(data_in[6]), .E(n293), .CP(clk), .Q(
        \input_value[7][6] ) );
  EDFQD1 \input_value_reg[7][5]  ( .D(data_in[5]), .E(n293), .CP(clk), .Q(
        \input_value[7][5] ) );
  EDFQD1 \input_value_reg[7][4]  ( .D(data_in[4]), .E(n293), .CP(clk), .Q(
        \input_value[7][4] ) );
  EDFQD1 \input_value_reg[7][3]  ( .D(data_in[3]), .E(n293), .CP(clk), .Q(
        \input_value[7][3] ) );
  EDFQD1 \input_value_reg[7][2]  ( .D(data_in[2]), .E(n293), .CP(clk), .Q(
        \input_value[7][2] ) );
  EDFQD1 \input_value_reg[7][1]  ( .D(data_in[1]), .E(n293), .CP(clk), .Q(
        \input_value[7][1] ) );
  EDFQD1 \input_value_reg[7][0]  ( .D(data_in[0]), .E(n293), .CP(clk), .Q(
        \input_value[7][0] ) );
  EDFQD1 \input_weight_reg[7][99]  ( .D(data_in[99]), .E(n422), .CP(clk), .Q(
        \input_weight[7][99] ) );
  EDFQD1 \input_weight_reg[7][100]  ( .D(data_in[100]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][100] ) );
  EDFQD1 \input_weight_reg[7][101]  ( .D(data_in[101]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][101] ) );
  EDFQD1 \input_weight_reg[7][102]  ( .D(data_in[102]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][102] ) );
  EDFQD1 \input_weight_reg[7][103]  ( .D(data_in[103]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][103] ) );
  EDFQD1 \input_weight_reg[7][104]  ( .D(data_in[104]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][104] ) );
  EDFQD1 \input_weight_reg[7][105]  ( .D(data_in[105]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][105] ) );
  EDFQD1 \input_weight_reg[7][106]  ( .D(data_in[106]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][106] ) );
  EDFQD1 \input_weight_reg[7][107]  ( .D(data_in[107]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][107] ) );
  EDFQD1 \input_weight_reg[7][108]  ( .D(data_in[108]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][108] ) );
  EDFQD1 \input_weight_reg[7][109]  ( .D(data_in[109]), .E(n422), .CP(clk), 
        .Q(\input_weight[7][109] ) );
  EDFQD1 \input_weight_reg[7][110]  ( .D(data_in[110]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][110] ) );
  EDFQD1 \input_weight_reg[7][111]  ( .D(data_in[111]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][111] ) );
  EDFQD1 \input_weight_reg[7][112]  ( .D(data_in[112]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][112] ) );
  EDFQD1 \input_weight_reg[7][113]  ( .D(data_in[113]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][113] ) );
  EDFQD1 \input_weight_reg[7][114]  ( .D(data_in[114]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][114] ) );
  EDFQD1 \input_weight_reg[7][115]  ( .D(data_in[115]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][115] ) );
  EDFQD1 \input_weight_reg[7][116]  ( .D(data_in[116]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][116] ) );
  EDFQD1 \input_weight_reg[7][117]  ( .D(data_in[117]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][117] ) );
  EDFQD1 \input_weight_reg[7][118]  ( .D(data_in[118]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][118] ) );
  EDFQD1 \input_weight_reg[7][119]  ( .D(data_in[119]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][119] ) );
  EDFQD1 \input_weight_reg[7][120]  ( .D(data_in[120]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][120] ) );
  EDFQD1 \input_weight_reg[7][121]  ( .D(data_in[121]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][121] ) );
  EDFQD1 \input_weight_reg[7][122]  ( .D(data_in[122]), .E(n421), .CP(clk), 
        .Q(\input_weight[7][122] ) );
  EDFQD1 \input_weight_reg[7][123]  ( .D(data_in[123]), .E(n420), .CP(clk), 
        .Q(\input_weight[7][123] ) );
  EDFQD1 \input_weight_reg[7][124]  ( .D(data_in[124]), .E(n420), .CP(clk), 
        .Q(\input_weight[7][124] ) );
  EDFQD1 \input_weight_reg[7][125]  ( .D(data_in[125]), .E(n420), .CP(clk), 
        .Q(\input_weight[7][125] ) );
  EDFQD1 \input_weight_reg[7][126]  ( .D(data_in[126]), .E(n420), .CP(clk), 
        .Q(\input_weight[7][126] ) );
  EDFQD1 \input_weight_reg[7][127]  ( .D(data_in[127]), .E(n420), .CP(clk), 
        .Q(\input_weight[7][127] ) );
  EDFQD1 \input_weight_reg[7][98]  ( .D(data_in[98]), .E(n420), .CP(clk), .Q(
        \input_weight[7][98] ) );
  EDFQD1 \input_weight_reg[7][97]  ( .D(data_in[97]), .E(n420), .CP(clk), .Q(
        \input_weight[7][97] ) );
  EDFQD1 \input_weight_reg[7][96]  ( .D(data_in[96]), .E(n420), .CP(clk), .Q(
        \input_weight[7][96] ) );
  EDFQD1 \input_weight_reg[7][95]  ( .D(data_in[95]), .E(n420), .CP(clk), .Q(
        \input_weight[7][95] ) );
  EDFQD1 \input_weight_reg[7][94]  ( .D(data_in[94]), .E(n420), .CP(clk), .Q(
        \input_weight[7][94] ) );
  EDFQD1 \input_weight_reg[7][93]  ( .D(data_in[93]), .E(n420), .CP(clk), .Q(
        \input_weight[7][93] ) );
  EDFQD1 \input_weight_reg[7][92]  ( .D(data_in[92]), .E(n420), .CP(clk), .Q(
        \input_weight[7][92] ) );
  EDFQD1 \input_weight_reg[7][91]  ( .D(data_in[91]), .E(n420), .CP(clk), .Q(
        \input_weight[7][91] ) );
  EDFQD1 \input_weight_reg[7][90]  ( .D(data_in[90]), .E(n419), .CP(clk), .Q(
        \input_weight[7][90] ) );
  EDFQD1 \input_weight_reg[7][89]  ( .D(data_in[89]), .E(n419), .CP(clk), .Q(
        \input_weight[7][89] ) );
  EDFQD1 \input_weight_reg[7][88]  ( .D(data_in[88]), .E(n419), .CP(clk), .Q(
        \input_weight[7][88] ) );
  EDFQD1 \input_weight_reg[7][87]  ( .D(data_in[87]), .E(n419), .CP(clk), .Q(
        \input_weight[7][87] ) );
  EDFQD1 \input_weight_reg[7][86]  ( .D(data_in[86]), .E(n419), .CP(clk), .Q(
        \input_weight[7][86] ) );
  EDFQD1 \input_weight_reg[7][85]  ( .D(data_in[85]), .E(n419), .CP(clk), .Q(
        \input_weight[7][85] ) );
  EDFQD1 \input_weight_reg[7][84]  ( .D(data_in[84]), .E(n419), .CP(clk), .Q(
        \input_weight[7][84] ) );
  EDFQD1 \input_weight_reg[7][83]  ( .D(data_in[83]), .E(n419), .CP(clk), .Q(
        \input_weight[7][83] ) );
  EDFQD1 \input_weight_reg[7][82]  ( .D(data_in[82]), .E(n419), .CP(clk), .Q(
        \input_weight[7][82] ) );
  EDFQD1 \input_weight_reg[7][81]  ( .D(data_in[81]), .E(n419), .CP(clk), .Q(
        \input_weight[7][81] ) );
  EDFQD1 \input_weight_reg[7][80]  ( .D(data_in[80]), .E(n419), .CP(clk), .Q(
        \input_weight[7][80] ) );
  EDFQD1 \input_weight_reg[7][79]  ( .D(data_in[79]), .E(n419), .CP(clk), .Q(
        \input_weight[7][79] ) );
  EDFQD1 \input_weight_reg[7][78]  ( .D(data_in[78]), .E(n419), .CP(clk), .Q(
        \input_weight[7][78] ) );
  EDFQD1 \input_weight_reg[7][77]  ( .D(data_in[77]), .E(n418), .CP(clk), .Q(
        \input_weight[7][77] ) );
  EDFQD1 \input_weight_reg[7][76]  ( .D(data_in[76]), .E(n418), .CP(clk), .Q(
        \input_weight[7][76] ) );
  EDFQD1 \input_weight_reg[7][75]  ( .D(data_in[75]), .E(n418), .CP(clk), .Q(
        \input_weight[7][75] ) );
  EDFQD1 \input_weight_reg[7][74]  ( .D(data_in[74]), .E(n418), .CP(clk), .Q(
        \input_weight[7][74] ) );
  EDFQD1 \input_weight_reg[7][73]  ( .D(data_in[73]), .E(n418), .CP(clk), .Q(
        \input_weight[7][73] ) );
  EDFQD1 \input_weight_reg[7][72]  ( .D(data_in[72]), .E(n418), .CP(clk), .Q(
        \input_weight[7][72] ) );
  EDFQD1 \input_weight_reg[7][71]  ( .D(data_in[71]), .E(n418), .CP(clk), .Q(
        \input_weight[7][71] ) );
  EDFQD1 \input_weight_reg[7][70]  ( .D(data_in[70]), .E(n418), .CP(clk), .Q(
        \input_weight[7][70] ) );
  EDFQD1 \input_weight_reg[7][69]  ( .D(data_in[69]), .E(n418), .CP(clk), .Q(
        \input_weight[7][69] ) );
  EDFQD1 \input_weight_reg[7][68]  ( .D(data_in[68]), .E(n418), .CP(clk), .Q(
        \input_weight[7][68] ) );
  EDFQD1 \input_weight_reg[7][67]  ( .D(data_in[67]), .E(n418), .CP(clk), .Q(
        \input_weight[7][67] ) );
  EDFQD1 \input_weight_reg[7][66]  ( .D(data_in[66]), .E(n418), .CP(clk), .Q(
        \input_weight[7][66] ) );
  EDFQD1 \input_weight_reg[7][65]  ( .D(data_in[65]), .E(n418), .CP(clk), .Q(
        \input_weight[7][65] ) );
  EDFQD1 \input_weight_reg[7][64]  ( .D(data_in[64]), .E(n417), .CP(clk), .Q(
        \input_weight[7][64] ) );
  EDFQD1 \input_weight_reg[7][63]  ( .D(data_in[63]), .E(n417), .CP(clk), .Q(
        \input_weight[7][63] ) );
  EDFQD1 \input_weight_reg[7][62]  ( .D(data_in[62]), .E(n417), .CP(clk), .Q(
        \input_weight[7][62] ) );
  EDFQD1 \input_weight_reg[7][61]  ( .D(data_in[61]), .E(n417), .CP(clk), .Q(
        \input_weight[7][61] ) );
  EDFQD1 \input_weight_reg[7][60]  ( .D(data_in[60]), .E(n417), .CP(clk), .Q(
        \input_weight[7][60] ) );
  EDFQD1 \input_weight_reg[7][59]  ( .D(data_in[59]), .E(n417), .CP(clk), .Q(
        \input_weight[7][59] ) );
  EDFQD1 \input_weight_reg[7][58]  ( .D(data_in[58]), .E(n417), .CP(clk), .Q(
        \input_weight[7][58] ) );
  EDFQD1 \input_weight_reg[7][57]  ( .D(data_in[57]), .E(n417), .CP(clk), .Q(
        \input_weight[7][57] ) );
  EDFQD1 \input_weight_reg[7][56]  ( .D(data_in[56]), .E(n417), .CP(clk), .Q(
        \input_weight[7][56] ) );
  EDFQD1 \input_weight_reg[7][55]  ( .D(data_in[55]), .E(n417), .CP(clk), .Q(
        \input_weight[7][55] ) );
  EDFQD1 \input_weight_reg[7][54]  ( .D(data_in[54]), .E(n417), .CP(clk), .Q(
        \input_weight[7][54] ) );
  EDFQD1 \input_weight_reg[7][53]  ( .D(data_in[53]), .E(n417), .CP(clk), .Q(
        \input_weight[7][53] ) );
  EDFQD1 \input_weight_reg[7][52]  ( .D(data_in[52]), .E(n417), .CP(clk), .Q(
        \input_weight[7][52] ) );
  EDFQD1 \input_weight_reg[7][51]  ( .D(data_in[51]), .E(n416), .CP(clk), .Q(
        \input_weight[7][51] ) );
  EDFQD1 \input_weight_reg[7][50]  ( .D(data_in[50]), .E(n416), .CP(clk), .Q(
        \input_weight[7][50] ) );
  EDFQD1 \input_weight_reg[7][49]  ( .D(data_in[49]), .E(n416), .CP(clk), .Q(
        \input_weight[7][49] ) );
  EDFQD1 \input_weight_reg[7][48]  ( .D(data_in[48]), .E(n416), .CP(clk), .Q(
        \input_weight[7][48] ) );
  EDFQD1 \input_weight_reg[7][47]  ( .D(data_in[47]), .E(n416), .CP(clk), .Q(
        \input_weight[7][47] ) );
  EDFQD1 \input_weight_reg[7][46]  ( .D(data_in[46]), .E(n416), .CP(clk), .Q(
        \input_weight[7][46] ) );
  EDFQD1 \input_weight_reg[7][45]  ( .D(data_in[45]), .E(n416), .CP(clk), .Q(
        \input_weight[7][45] ) );
  EDFQD1 \input_weight_reg[7][44]  ( .D(data_in[44]), .E(n416), .CP(clk), .Q(
        \input_weight[7][44] ) );
  EDFQD1 \input_weight_reg[7][43]  ( .D(data_in[43]), .E(n416), .CP(clk), .Q(
        \input_weight[7][43] ) );
  EDFQD1 \input_weight_reg[7][42]  ( .D(data_in[42]), .E(n416), .CP(clk), .Q(
        \input_weight[7][42] ) );
  EDFQD1 \input_weight_reg[7][41]  ( .D(data_in[41]), .E(n416), .CP(clk), .Q(
        \input_weight[7][41] ) );
  EDFQD1 \input_weight_reg[7][40]  ( .D(data_in[40]), .E(n416), .CP(clk), .Q(
        \input_weight[7][40] ) );
  EDFQD1 \input_weight_reg[7][39]  ( .D(data_in[39]), .E(n416), .CP(clk), .Q(
        \input_weight[7][39] ) );
  EDFQD1 \input_weight_reg[7][38]  ( .D(data_in[38]), .E(n415), .CP(clk), .Q(
        \input_weight[7][38] ) );
  EDFQD1 \input_weight_reg[7][37]  ( .D(data_in[37]), .E(n415), .CP(clk), .Q(
        \input_weight[7][37] ) );
  EDFQD1 \input_weight_reg[7][36]  ( .D(data_in[36]), .E(n415), .CP(clk), .Q(
        \input_weight[7][36] ) );
  EDFQD1 \input_weight_reg[7][35]  ( .D(data_in[35]), .E(n415), .CP(clk), .Q(
        \input_weight[7][35] ) );
  EDFQD1 \input_weight_reg[7][34]  ( .D(data_in[34]), .E(n415), .CP(clk), .Q(
        \input_weight[7][34] ) );
  EDFQD1 \input_weight_reg[7][33]  ( .D(data_in[33]), .E(n415), .CP(clk), .Q(
        \input_weight[7][33] ) );
  EDFQD1 \input_weight_reg[7][32]  ( .D(data_in[32]), .E(n415), .CP(clk), .Q(
        \input_weight[7][32] ) );
  EDFQD1 \input_weight_reg[7][31]  ( .D(data_in[31]), .E(n415), .CP(clk), .Q(
        \input_weight[7][31] ) );
  EDFQD1 \input_weight_reg[7][30]  ( .D(data_in[30]), .E(n415), .CP(clk), .Q(
        \input_weight[7][30] ) );
  EDFQD1 \input_weight_reg[7][29]  ( .D(data_in[29]), .E(n415), .CP(clk), .Q(
        \input_weight[7][29] ) );
  EDFQD1 \input_weight_reg[7][28]  ( .D(data_in[28]), .E(n415), .CP(clk), .Q(
        \input_weight[7][28] ) );
  EDFQD1 \input_weight_reg[7][27]  ( .D(data_in[27]), .E(n415), .CP(clk), .Q(
        \input_weight[7][27] ) );
  EDFQD1 \input_weight_reg[7][26]  ( .D(data_in[26]), .E(n415), .CP(clk), .Q(
        \input_weight[7][26] ) );
  EDFQD1 \input_weight_reg[7][25]  ( .D(data_in[25]), .E(n414), .CP(clk), .Q(
        \input_weight[7][25] ) );
  EDFQD1 \input_weight_reg[7][24]  ( .D(data_in[24]), .E(n414), .CP(clk), .Q(
        \input_weight[7][24] ) );
  EDFQD1 \input_weight_reg[7][23]  ( .D(data_in[23]), .E(n414), .CP(clk), .Q(
        \input_weight[7][23] ) );
  EDFQD1 \input_weight_reg[7][22]  ( .D(data_in[22]), .E(n414), .CP(clk), .Q(
        \input_weight[7][22] ) );
  EDFQD1 \input_weight_reg[7][21]  ( .D(data_in[21]), .E(n414), .CP(clk), .Q(
        \input_weight[7][21] ) );
  EDFQD1 \input_weight_reg[7][20]  ( .D(data_in[20]), .E(n414), .CP(clk), .Q(
        \input_weight[7][20] ) );
  EDFQD1 \input_weight_reg[7][19]  ( .D(data_in[19]), .E(n414), .CP(clk), .Q(
        \input_weight[7][19] ) );
  EDFQD1 \input_weight_reg[7][18]  ( .D(data_in[18]), .E(n414), .CP(clk), .Q(
        \input_weight[7][18] ) );
  EDFQD1 \input_weight_reg[7][17]  ( .D(data_in[17]), .E(n414), .CP(clk), .Q(
        \input_weight[7][17] ) );
  EDFQD1 \input_weight_reg[7][16]  ( .D(data_in[16]), .E(n414), .CP(clk), .Q(
        \input_weight[7][16] ) );
  EDFQD1 \input_weight_reg[7][15]  ( .D(data_in[15]), .E(n414), .CP(clk), .Q(
        \input_weight[7][15] ) );
  EDFQD1 \input_weight_reg[7][14]  ( .D(data_in[14]), .E(n414), .CP(clk), .Q(
        \input_weight[7][14] ) );
  EDFQD1 \input_weight_reg[7][13]  ( .D(data_in[13]), .E(n414), .CP(clk), .Q(
        \input_weight[7][13] ) );
  EDFQD1 \input_weight_reg[7][12]  ( .D(data_in[12]), .E(n413), .CP(clk), .Q(
        \input_weight[7][12] ) );
  EDFQD1 \input_weight_reg[7][11]  ( .D(data_in[11]), .E(n413), .CP(clk), .Q(
        \input_weight[7][11] ) );
  EDFQD1 \input_weight_reg[7][10]  ( .D(data_in[10]), .E(n413), .CP(clk), .Q(
        \input_weight[7][10] ) );
  EDFQD1 \input_weight_reg[7][9]  ( .D(data_in[9]), .E(n413), .CP(clk), .Q(
        \input_weight[7][9] ) );
  EDFQD1 \input_weight_reg[7][8]  ( .D(data_in[8]), .E(n413), .CP(clk), .Q(
        \input_weight[7][8] ) );
  EDFQD1 \input_weight_reg[7][7]  ( .D(data_in[7]), .E(n413), .CP(clk), .Q(
        \input_weight[7][7] ) );
  EDFQD1 \input_weight_reg[7][6]  ( .D(data_in[6]), .E(n413), .CP(clk), .Q(
        \input_weight[7][6] ) );
  EDFQD1 \input_weight_reg[7][5]  ( .D(data_in[5]), .E(n413), .CP(clk), .Q(
        \input_weight[7][5] ) );
  EDFQD1 \input_weight_reg[7][4]  ( .D(data_in[4]), .E(n413), .CP(clk), .Q(
        \input_weight[7][4] ) );
  EDFQD1 \input_weight_reg[7][3]  ( .D(data_in[3]), .E(n413), .CP(clk), .Q(
        \input_weight[7][3] ) );
  EDFQD1 \input_weight_reg[7][2]  ( .D(data_in[2]), .E(n413), .CP(clk), .Q(
        \input_weight[7][2] ) );
  EDFQD1 \input_weight_reg[7][1]  ( .D(data_in[1]), .E(n413), .CP(clk), .Q(
        \input_weight[7][1] ) );
  EDFQD1 \input_weight_reg[7][0]  ( .D(data_in[0]), .E(n413), .CP(clk), .Q(
        \input_weight[7][0] ) );
  EDFQD1 \input_value_reg[5][99]  ( .D(data_in[99]), .E(n332), .CP(clk), .Q(
        \input_value[5][99] ) );
  EDFQD1 \input_value_reg[5][100]  ( .D(data_in[100]), .E(n332), .CP(clk), .Q(
        \input_value[5][100] ) );
  EDFQD1 \input_value_reg[5][101]  ( .D(data_in[101]), .E(n332), .CP(clk), .Q(
        \input_value[5][101] ) );
  EDFQD1 \input_value_reg[5][102]  ( .D(data_in[102]), .E(n332), .CP(clk), .Q(
        \input_value[5][102] ) );
  EDFQD1 \input_value_reg[5][103]  ( .D(data_in[103]), .E(n332), .CP(clk), .Q(
        \input_value[5][103] ) );
  EDFQD1 \input_value_reg[5][104]  ( .D(data_in[104]), .E(n332), .CP(clk), .Q(
        \input_value[5][104] ) );
  EDFQD1 \input_value_reg[5][105]  ( .D(data_in[105]), .E(n332), .CP(clk), .Q(
        \input_value[5][105] ) );
  EDFQD1 \input_value_reg[5][106]  ( .D(data_in[106]), .E(n332), .CP(clk), .Q(
        \input_value[5][106] ) );
  EDFQD1 \input_value_reg[5][107]  ( .D(data_in[107]), .E(n332), .CP(clk), .Q(
        \input_value[5][107] ) );
  EDFQD1 \input_value_reg[5][108]  ( .D(data_in[108]), .E(n332), .CP(clk), .Q(
        \input_value[5][108] ) );
  EDFQD1 \input_value_reg[5][109]  ( .D(data_in[109]), .E(n332), .CP(clk), .Q(
        \input_value[5][109] ) );
  EDFQD1 \input_value_reg[5][110]  ( .D(data_in[110]), .E(n331), .CP(clk), .Q(
        \input_value[5][110] ) );
  EDFQD1 \input_value_reg[5][111]  ( .D(data_in[111]), .E(n331), .CP(clk), .Q(
        \input_value[5][111] ) );
  EDFQD1 \input_value_reg[5][112]  ( .D(data_in[112]), .E(n331), .CP(clk), .Q(
        \input_value[5][112] ) );
  EDFQD1 \input_value_reg[5][113]  ( .D(data_in[113]), .E(n331), .CP(clk), .Q(
        \input_value[5][113] ) );
  EDFQD1 \input_value_reg[5][114]  ( .D(data_in[114]), .E(n331), .CP(clk), .Q(
        \input_value[5][114] ) );
  EDFQD1 \input_value_reg[5][115]  ( .D(data_in[115]), .E(n331), .CP(clk), .Q(
        \input_value[5][115] ) );
  EDFQD1 \input_value_reg[5][116]  ( .D(data_in[116]), .E(n331), .CP(clk), .Q(
        \input_value[5][116] ) );
  EDFQD1 \input_value_reg[5][117]  ( .D(data_in[117]), .E(n331), .CP(clk), .Q(
        \input_value[5][117] ) );
  EDFQD1 \input_value_reg[5][118]  ( .D(data_in[118]), .E(n331), .CP(clk), .Q(
        \input_value[5][118] ) );
  EDFQD1 \input_value_reg[5][119]  ( .D(data_in[119]), .E(n331), .CP(clk), .Q(
        \input_value[5][119] ) );
  EDFQD1 \input_value_reg[5][120]  ( .D(data_in[120]), .E(n331), .CP(clk), .Q(
        \input_value[5][120] ) );
  EDFQD1 \input_value_reg[5][121]  ( .D(data_in[121]), .E(n331), .CP(clk), .Q(
        \input_value[5][121] ) );
  EDFQD1 \input_value_reg[5][122]  ( .D(data_in[122]), .E(n331), .CP(clk), .Q(
        \input_value[5][122] ) );
  EDFQD1 \input_value_reg[5][123]  ( .D(data_in[123]), .E(n330), .CP(clk), .Q(
        \input_value[5][123] ) );
  EDFQD1 \input_value_reg[5][124]  ( .D(data_in[124]), .E(n330), .CP(clk), .Q(
        \input_value[5][124] ) );
  EDFQD1 \input_value_reg[5][125]  ( .D(data_in[125]), .E(n330), .CP(clk), .Q(
        \input_value[5][125] ) );
  EDFQD1 \input_value_reg[5][126]  ( .D(data_in[126]), .E(n330), .CP(clk), .Q(
        \input_value[5][126] ) );
  EDFQD1 \input_value_reg[5][127]  ( .D(data_in[127]), .E(n330), .CP(clk), .Q(
        \input_value[5][127] ) );
  EDFQD1 \input_value_reg[5][98]  ( .D(data_in[98]), .E(n330), .CP(clk), .Q(
        \input_value[5][98] ) );
  EDFQD1 \input_value_reg[5][97]  ( .D(data_in[97]), .E(n330), .CP(clk), .Q(
        \input_value[5][97] ) );
  EDFQD1 \input_value_reg[5][96]  ( .D(data_in[96]), .E(n330), .CP(clk), .Q(
        \input_value[5][96] ) );
  EDFQD1 \input_value_reg[5][95]  ( .D(data_in[95]), .E(n330), .CP(clk), .Q(
        \input_value[5][95] ) );
  EDFQD1 \input_value_reg[5][94]  ( .D(data_in[94]), .E(n330), .CP(clk), .Q(
        \input_value[5][94] ) );
  EDFQD1 \input_value_reg[5][93]  ( .D(data_in[93]), .E(n330), .CP(clk), .Q(
        \input_value[5][93] ) );
  EDFQD1 \input_value_reg[5][92]  ( .D(data_in[92]), .E(n330), .CP(clk), .Q(
        \input_value[5][92] ) );
  EDFQD1 \input_value_reg[5][91]  ( .D(data_in[91]), .E(n330), .CP(clk), .Q(
        \input_value[5][91] ) );
  EDFQD1 \input_value_reg[5][90]  ( .D(data_in[90]), .E(n329), .CP(clk), .Q(
        \input_value[5][90] ) );
  EDFQD1 \input_value_reg[5][89]  ( .D(data_in[89]), .E(n329), .CP(clk), .Q(
        \input_value[5][89] ) );
  EDFQD1 \input_value_reg[5][88]  ( .D(data_in[88]), .E(n329), .CP(clk), .Q(
        \input_value[5][88] ) );
  EDFQD1 \input_value_reg[5][87]  ( .D(data_in[87]), .E(n329), .CP(clk), .Q(
        \input_value[5][87] ) );
  EDFQD1 \input_value_reg[5][86]  ( .D(data_in[86]), .E(n329), .CP(clk), .Q(
        \input_value[5][86] ) );
  EDFQD1 \input_value_reg[5][85]  ( .D(data_in[85]), .E(n329), .CP(clk), .Q(
        \input_value[5][85] ) );
  EDFQD1 \input_value_reg[5][84]  ( .D(data_in[84]), .E(n329), .CP(clk), .Q(
        \input_value[5][84] ) );
  EDFQD1 \input_value_reg[5][83]  ( .D(data_in[83]), .E(n329), .CP(clk), .Q(
        \input_value[5][83] ) );
  EDFQD1 \input_value_reg[5][82]  ( .D(data_in[82]), .E(n329), .CP(clk), .Q(
        \input_value[5][82] ) );
  EDFQD1 \input_value_reg[5][81]  ( .D(data_in[81]), .E(n329), .CP(clk), .Q(
        \input_value[5][81] ) );
  EDFQD1 \input_value_reg[5][80]  ( .D(data_in[80]), .E(n329), .CP(clk), .Q(
        \input_value[5][80] ) );
  EDFQD1 \input_value_reg[5][79]  ( .D(data_in[79]), .E(n329), .CP(clk), .Q(
        \input_value[5][79] ) );
  EDFQD1 \input_value_reg[5][78]  ( .D(data_in[78]), .E(n329), .CP(clk), .Q(
        \input_value[5][78] ) );
  EDFQD1 \input_value_reg[5][77]  ( .D(data_in[77]), .E(n328), .CP(clk), .Q(
        \input_value[5][77] ) );
  EDFQD1 \input_value_reg[5][76]  ( .D(data_in[76]), .E(n328), .CP(clk), .Q(
        \input_value[5][76] ) );
  EDFQD1 \input_value_reg[5][75]  ( .D(data_in[75]), .E(n328), .CP(clk), .Q(
        \input_value[5][75] ) );
  EDFQD1 \input_value_reg[5][74]  ( .D(data_in[74]), .E(n328), .CP(clk), .Q(
        \input_value[5][74] ) );
  EDFQD1 \input_value_reg[5][73]  ( .D(data_in[73]), .E(n328), .CP(clk), .Q(
        \input_value[5][73] ) );
  EDFQD1 \input_value_reg[5][72]  ( .D(data_in[72]), .E(n328), .CP(clk), .Q(
        \input_value[5][72] ) );
  EDFQD1 \input_value_reg[5][71]  ( .D(data_in[71]), .E(n328), .CP(clk), .Q(
        \input_value[5][71] ) );
  EDFQD1 \input_value_reg[5][70]  ( .D(data_in[70]), .E(n328), .CP(clk), .Q(
        \input_value[5][70] ) );
  EDFQD1 \input_value_reg[5][69]  ( .D(data_in[69]), .E(n328), .CP(clk), .Q(
        \input_value[5][69] ) );
  EDFQD1 \input_value_reg[5][68]  ( .D(data_in[68]), .E(n328), .CP(clk), .Q(
        \input_value[5][68] ) );
  EDFQD1 \input_value_reg[5][67]  ( .D(data_in[67]), .E(n328), .CP(clk), .Q(
        \input_value[5][67] ) );
  EDFQD1 \input_value_reg[5][66]  ( .D(data_in[66]), .E(n328), .CP(clk), .Q(
        \input_value[5][66] ) );
  EDFQD1 \input_value_reg[5][65]  ( .D(data_in[65]), .E(n328), .CP(clk), .Q(
        \input_value[5][65] ) );
  EDFQD1 \input_value_reg[5][64]  ( .D(data_in[64]), .E(n327), .CP(clk), .Q(
        \input_value[5][64] ) );
  EDFQD1 \input_value_reg[5][63]  ( .D(data_in[63]), .E(n327), .CP(clk), .Q(
        \input_value[5][63] ) );
  EDFQD1 \input_value_reg[5][62]  ( .D(data_in[62]), .E(n327), .CP(clk), .Q(
        \input_value[5][62] ) );
  EDFQD1 \input_value_reg[5][61]  ( .D(data_in[61]), .E(n327), .CP(clk), .Q(
        \input_value[5][61] ) );
  EDFQD1 \input_value_reg[5][60]  ( .D(data_in[60]), .E(n327), .CP(clk), .Q(
        \input_value[5][60] ) );
  EDFQD1 \input_value_reg[5][59]  ( .D(data_in[59]), .E(n327), .CP(clk), .Q(
        \input_value[5][59] ) );
  EDFQD1 \input_value_reg[5][58]  ( .D(data_in[58]), .E(n327), .CP(clk), .Q(
        \input_value[5][58] ) );
  EDFQD1 \input_value_reg[5][57]  ( .D(data_in[57]), .E(n327), .CP(clk), .Q(
        \input_value[5][57] ) );
  EDFQD1 \input_value_reg[5][56]  ( .D(data_in[56]), .E(n327), .CP(clk), .Q(
        \input_value[5][56] ) );
  EDFQD1 \input_value_reg[5][55]  ( .D(data_in[55]), .E(n327), .CP(clk), .Q(
        \input_value[5][55] ) );
  EDFQD1 \input_value_reg[5][54]  ( .D(data_in[54]), .E(n327), .CP(clk), .Q(
        \input_value[5][54] ) );
  EDFQD1 \input_value_reg[5][53]  ( .D(data_in[53]), .E(n327), .CP(clk), .Q(
        \input_value[5][53] ) );
  EDFQD1 \input_value_reg[5][52]  ( .D(data_in[52]), .E(n327), .CP(clk), .Q(
        \input_value[5][52] ) );
  EDFQD1 \input_value_reg[5][51]  ( .D(data_in[51]), .E(n326), .CP(clk), .Q(
        \input_value[5][51] ) );
  EDFQD1 \input_value_reg[5][50]  ( .D(data_in[50]), .E(n326), .CP(clk), .Q(
        \input_value[5][50] ) );
  EDFQD1 \input_value_reg[5][49]  ( .D(data_in[49]), .E(n326), .CP(clk), .Q(
        \input_value[5][49] ) );
  EDFQD1 \input_value_reg[5][48]  ( .D(data_in[48]), .E(n326), .CP(clk), .Q(
        \input_value[5][48] ) );
  EDFQD1 \input_value_reg[5][47]  ( .D(data_in[47]), .E(n326), .CP(clk), .Q(
        \input_value[5][47] ) );
  EDFQD1 \input_value_reg[5][46]  ( .D(data_in[46]), .E(n326), .CP(clk), .Q(
        \input_value[5][46] ) );
  EDFQD1 \input_value_reg[5][45]  ( .D(data_in[45]), .E(n326), .CP(clk), .Q(
        \input_value[5][45] ) );
  EDFQD1 \input_value_reg[5][44]  ( .D(data_in[44]), .E(n326), .CP(clk), .Q(
        \input_value[5][44] ) );
  EDFQD1 \input_value_reg[5][43]  ( .D(data_in[43]), .E(n326), .CP(clk), .Q(
        \input_value[5][43] ) );
  EDFQD1 \input_value_reg[5][42]  ( .D(data_in[42]), .E(n326), .CP(clk), .Q(
        \input_value[5][42] ) );
  EDFQD1 \input_value_reg[5][41]  ( .D(data_in[41]), .E(n326), .CP(clk), .Q(
        \input_value[5][41] ) );
  EDFQD1 \input_value_reg[5][40]  ( .D(data_in[40]), .E(n326), .CP(clk), .Q(
        \input_value[5][40] ) );
  EDFQD1 \input_value_reg[5][39]  ( .D(data_in[39]), .E(n326), .CP(clk), .Q(
        \input_value[5][39] ) );
  EDFQD1 \input_value_reg[5][38]  ( .D(data_in[38]), .E(n325), .CP(clk), .Q(
        \input_value[5][38] ) );
  EDFQD1 \input_value_reg[5][37]  ( .D(data_in[37]), .E(n325), .CP(clk), .Q(
        \input_value[5][37] ) );
  EDFQD1 \input_value_reg[5][36]  ( .D(data_in[36]), .E(n325), .CP(clk), .Q(
        \input_value[5][36] ) );
  EDFQD1 \input_value_reg[5][35]  ( .D(data_in[35]), .E(n325), .CP(clk), .Q(
        \input_value[5][35] ) );
  EDFQD1 \input_value_reg[5][34]  ( .D(data_in[34]), .E(n325), .CP(clk), .Q(
        \input_value[5][34] ) );
  EDFQD1 \input_value_reg[5][33]  ( .D(data_in[33]), .E(n325), .CP(clk), .Q(
        \input_value[5][33] ) );
  EDFQD1 \input_value_reg[5][32]  ( .D(data_in[32]), .E(n325), .CP(clk), .Q(
        \input_value[5][32] ) );
  EDFQD1 \input_value_reg[5][31]  ( .D(data_in[31]), .E(n325), .CP(clk), .Q(
        \input_value[5][31] ) );
  EDFQD1 \input_value_reg[5][30]  ( .D(data_in[30]), .E(n325), .CP(clk), .Q(
        \input_value[5][30] ) );
  EDFQD1 \input_value_reg[5][29]  ( .D(data_in[29]), .E(n325), .CP(clk), .Q(
        \input_value[5][29] ) );
  EDFQD1 \input_value_reg[5][28]  ( .D(data_in[28]), .E(n325), .CP(clk), .Q(
        \input_value[5][28] ) );
  EDFQD1 \input_value_reg[5][27]  ( .D(data_in[27]), .E(n325), .CP(clk), .Q(
        \input_value[5][27] ) );
  EDFQD1 \input_value_reg[5][26]  ( .D(data_in[26]), .E(n325), .CP(clk), .Q(
        \input_value[5][26] ) );
  EDFQD1 \input_value_reg[5][25]  ( .D(data_in[25]), .E(n324), .CP(clk), .Q(
        \input_value[5][25] ) );
  EDFQD1 \input_value_reg[5][24]  ( .D(data_in[24]), .E(n324), .CP(clk), .Q(
        \input_value[5][24] ) );
  EDFQD1 \input_value_reg[5][23]  ( .D(data_in[23]), .E(n324), .CP(clk), .Q(
        \input_value[5][23] ) );
  EDFQD1 \input_value_reg[5][22]  ( .D(data_in[22]), .E(n324), .CP(clk), .Q(
        \input_value[5][22] ) );
  EDFQD1 \input_value_reg[5][21]  ( .D(data_in[21]), .E(n324), .CP(clk), .Q(
        \input_value[5][21] ) );
  EDFQD1 \input_value_reg[5][20]  ( .D(data_in[20]), .E(n324), .CP(clk), .Q(
        \input_value[5][20] ) );
  EDFQD1 \input_value_reg[5][19]  ( .D(data_in[19]), .E(n324), .CP(clk), .Q(
        \input_value[5][19] ) );
  EDFQD1 \input_value_reg[5][18]  ( .D(data_in[18]), .E(n324), .CP(clk), .Q(
        \input_value[5][18] ) );
  EDFQD1 \input_value_reg[5][17]  ( .D(data_in[17]), .E(n324), .CP(clk), .Q(
        \input_value[5][17] ) );
  EDFQD1 \input_value_reg[5][16]  ( .D(data_in[16]), .E(n324), .CP(clk), .Q(
        \input_value[5][16] ) );
  EDFQD1 \input_value_reg[5][15]  ( .D(data_in[15]), .E(n324), .CP(clk), .Q(
        \input_value[5][15] ) );
  EDFQD1 \input_value_reg[5][14]  ( .D(data_in[14]), .E(n324), .CP(clk), .Q(
        \input_value[5][14] ) );
  EDFQD1 \input_value_reg[5][13]  ( .D(data_in[13]), .E(n324), .CP(clk), .Q(
        \input_value[5][13] ) );
  EDFQD1 \input_value_reg[5][12]  ( .D(data_in[12]), .E(n323), .CP(clk), .Q(
        \input_value[5][12] ) );
  EDFQD1 \input_value_reg[5][11]  ( .D(data_in[11]), .E(n323), .CP(clk), .Q(
        \input_value[5][11] ) );
  EDFQD1 \input_value_reg[5][10]  ( .D(data_in[10]), .E(n323), .CP(clk), .Q(
        \input_value[5][10] ) );
  EDFQD1 \input_value_reg[5][9]  ( .D(data_in[9]), .E(n323), .CP(clk), .Q(
        \input_value[5][9] ) );
  EDFQD1 \input_value_reg[5][8]  ( .D(data_in[8]), .E(n323), .CP(clk), .Q(
        \input_value[5][8] ) );
  EDFQD1 \input_value_reg[5][7]  ( .D(data_in[7]), .E(n323), .CP(clk), .Q(
        \input_value[5][7] ) );
  EDFQD1 \input_value_reg[5][6]  ( .D(data_in[6]), .E(n323), .CP(clk), .Q(
        \input_value[5][6] ) );
  EDFQD1 \input_value_reg[5][5]  ( .D(data_in[5]), .E(n323), .CP(clk), .Q(
        \input_value[5][5] ) );
  EDFQD1 \input_value_reg[5][4]  ( .D(data_in[4]), .E(n323), .CP(clk), .Q(
        \input_value[5][4] ) );
  EDFQD1 \input_value_reg[5][3]  ( .D(data_in[3]), .E(n323), .CP(clk), .Q(
        \input_value[5][3] ) );
  EDFQD1 \input_value_reg[5][2]  ( .D(data_in[2]), .E(n323), .CP(clk), .Q(
        \input_value[5][2] ) );
  EDFQD1 \input_value_reg[5][1]  ( .D(data_in[1]), .E(n323), .CP(clk), .Q(
        \input_value[5][1] ) );
  EDFQD1 \input_value_reg[5][0]  ( .D(data_in[0]), .E(n323), .CP(clk), .Q(
        \input_value[5][0] ) );
  EDFQD1 \input_weight_reg[5][99]  ( .D(data_in[99]), .E(n452), .CP(clk), .Q(
        \input_weight[5][99] ) );
  EDFQD1 \input_weight_reg[5][100]  ( .D(data_in[100]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][100] ) );
  EDFQD1 \input_weight_reg[5][101]  ( .D(data_in[101]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][101] ) );
  EDFQD1 \input_weight_reg[5][102]  ( .D(data_in[102]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][102] ) );
  EDFQD1 \input_weight_reg[5][103]  ( .D(data_in[103]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][103] ) );
  EDFQD1 \input_weight_reg[5][104]  ( .D(data_in[104]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][104] ) );
  EDFQD1 \input_weight_reg[5][105]  ( .D(data_in[105]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][105] ) );
  EDFQD1 \input_weight_reg[5][106]  ( .D(data_in[106]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][106] ) );
  EDFQD1 \input_weight_reg[5][107]  ( .D(data_in[107]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][107] ) );
  EDFQD1 \input_weight_reg[5][108]  ( .D(data_in[108]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][108] ) );
  EDFQD1 \input_weight_reg[5][109]  ( .D(data_in[109]), .E(n452), .CP(clk), 
        .Q(\input_weight[5][109] ) );
  EDFQD1 \input_weight_reg[5][110]  ( .D(data_in[110]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][110] ) );
  EDFQD1 \input_weight_reg[5][111]  ( .D(data_in[111]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][111] ) );
  EDFQD1 \input_weight_reg[5][112]  ( .D(data_in[112]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][112] ) );
  EDFQD1 \input_weight_reg[5][113]  ( .D(data_in[113]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][113] ) );
  EDFQD1 \input_weight_reg[5][114]  ( .D(data_in[114]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][114] ) );
  EDFQD1 \input_weight_reg[5][115]  ( .D(data_in[115]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][115] ) );
  EDFQD1 \input_weight_reg[5][116]  ( .D(data_in[116]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][116] ) );
  EDFQD1 \input_weight_reg[5][117]  ( .D(data_in[117]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][117] ) );
  EDFQD1 \input_weight_reg[5][118]  ( .D(data_in[118]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][118] ) );
  EDFQD1 \input_weight_reg[5][119]  ( .D(data_in[119]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][119] ) );
  EDFQD1 \input_weight_reg[5][120]  ( .D(data_in[120]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][120] ) );
  EDFQD1 \input_weight_reg[5][121]  ( .D(data_in[121]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][121] ) );
  EDFQD1 \input_weight_reg[5][122]  ( .D(data_in[122]), .E(n451), .CP(clk), 
        .Q(\input_weight[5][122] ) );
  EDFQD1 \input_weight_reg[5][123]  ( .D(data_in[123]), .E(n450), .CP(clk), 
        .Q(\input_weight[5][123] ) );
  EDFQD1 \input_weight_reg[5][124]  ( .D(data_in[124]), .E(n450), .CP(clk), 
        .Q(\input_weight[5][124] ) );
  EDFQD1 \input_weight_reg[5][125]  ( .D(data_in[125]), .E(n450), .CP(clk), 
        .Q(\input_weight[5][125] ) );
  EDFQD1 \input_weight_reg[5][126]  ( .D(data_in[126]), .E(n450), .CP(clk), 
        .Q(\input_weight[5][126] ) );
  EDFQD1 \input_weight_reg[5][127]  ( .D(data_in[127]), .E(n450), .CP(clk), 
        .Q(\input_weight[5][127] ) );
  EDFQD1 \input_weight_reg[5][98]  ( .D(data_in[98]), .E(n450), .CP(clk), .Q(
        \input_weight[5][98] ) );
  EDFQD1 \input_weight_reg[5][97]  ( .D(data_in[97]), .E(n450), .CP(clk), .Q(
        \input_weight[5][97] ) );
  EDFQD1 \input_weight_reg[5][96]  ( .D(data_in[96]), .E(n450), .CP(clk), .Q(
        \input_weight[5][96] ) );
  EDFQD1 \input_weight_reg[5][95]  ( .D(data_in[95]), .E(n450), .CP(clk), .Q(
        \input_weight[5][95] ) );
  EDFQD1 \input_weight_reg[5][94]  ( .D(data_in[94]), .E(n450), .CP(clk), .Q(
        \input_weight[5][94] ) );
  EDFQD1 \input_weight_reg[5][93]  ( .D(data_in[93]), .E(n450), .CP(clk), .Q(
        \input_weight[5][93] ) );
  EDFQD1 \input_weight_reg[5][92]  ( .D(data_in[92]), .E(n450), .CP(clk), .Q(
        \input_weight[5][92] ) );
  EDFQD1 \input_weight_reg[5][91]  ( .D(data_in[91]), .E(n450), .CP(clk), .Q(
        \input_weight[5][91] ) );
  EDFQD1 \input_weight_reg[5][90]  ( .D(data_in[90]), .E(n449), .CP(clk), .Q(
        \input_weight[5][90] ) );
  EDFQD1 \input_weight_reg[5][89]  ( .D(data_in[89]), .E(n449), .CP(clk), .Q(
        \input_weight[5][89] ) );
  EDFQD1 \input_weight_reg[5][88]  ( .D(data_in[88]), .E(n449), .CP(clk), .Q(
        \input_weight[5][88] ) );
  EDFQD1 \input_weight_reg[5][87]  ( .D(data_in[87]), .E(n449), .CP(clk), .Q(
        \input_weight[5][87] ) );
  EDFQD1 \input_weight_reg[5][86]  ( .D(data_in[86]), .E(n449), .CP(clk), .Q(
        \input_weight[5][86] ) );
  EDFQD1 \input_weight_reg[5][85]  ( .D(data_in[85]), .E(n449), .CP(clk), .Q(
        \input_weight[5][85] ) );
  EDFQD1 \input_weight_reg[5][84]  ( .D(data_in[84]), .E(n449), .CP(clk), .Q(
        \input_weight[5][84] ) );
  EDFQD1 \input_weight_reg[5][83]  ( .D(data_in[83]), .E(n449), .CP(clk), .Q(
        \input_weight[5][83] ) );
  EDFQD1 \input_weight_reg[5][82]  ( .D(data_in[82]), .E(n449), .CP(clk), .Q(
        \input_weight[5][82] ) );
  EDFQD1 \input_weight_reg[5][81]  ( .D(data_in[81]), .E(n449), .CP(clk), .Q(
        \input_weight[5][81] ) );
  EDFQD1 \input_weight_reg[5][80]  ( .D(data_in[80]), .E(n449), .CP(clk), .Q(
        \input_weight[5][80] ) );
  EDFQD1 \input_weight_reg[5][79]  ( .D(data_in[79]), .E(n449), .CP(clk), .Q(
        \input_weight[5][79] ) );
  EDFQD1 \input_weight_reg[5][78]  ( .D(data_in[78]), .E(n449), .CP(clk), .Q(
        \input_weight[5][78] ) );
  EDFQD1 \input_weight_reg[5][77]  ( .D(data_in[77]), .E(n448), .CP(clk), .Q(
        \input_weight[5][77] ) );
  EDFQD1 \input_weight_reg[5][76]  ( .D(data_in[76]), .E(n448), .CP(clk), .Q(
        \input_weight[5][76] ) );
  EDFQD1 \input_weight_reg[5][75]  ( .D(data_in[75]), .E(n448), .CP(clk), .Q(
        \input_weight[5][75] ) );
  EDFQD1 \input_weight_reg[5][74]  ( .D(data_in[74]), .E(n448), .CP(clk), .Q(
        \input_weight[5][74] ) );
  EDFQD1 \input_weight_reg[5][73]  ( .D(data_in[73]), .E(n448), .CP(clk), .Q(
        \input_weight[5][73] ) );
  EDFQD1 \input_weight_reg[5][72]  ( .D(data_in[72]), .E(n448), .CP(clk), .Q(
        \input_weight[5][72] ) );
  EDFQD1 \input_weight_reg[5][71]  ( .D(data_in[71]), .E(n448), .CP(clk), .Q(
        \input_weight[5][71] ) );
  EDFQD1 \input_weight_reg[5][70]  ( .D(data_in[70]), .E(n448), .CP(clk), .Q(
        \input_weight[5][70] ) );
  EDFQD1 \input_weight_reg[5][69]  ( .D(data_in[69]), .E(n448), .CP(clk), .Q(
        \input_weight[5][69] ) );
  EDFQD1 \input_weight_reg[5][68]  ( .D(data_in[68]), .E(n448), .CP(clk), .Q(
        \input_weight[5][68] ) );
  EDFQD1 \input_weight_reg[5][67]  ( .D(data_in[67]), .E(n448), .CP(clk), .Q(
        \input_weight[5][67] ) );
  EDFQD1 \input_weight_reg[5][66]  ( .D(data_in[66]), .E(n448), .CP(clk), .Q(
        \input_weight[5][66] ) );
  EDFQD1 \input_weight_reg[5][65]  ( .D(data_in[65]), .E(n448), .CP(clk), .Q(
        \input_weight[5][65] ) );
  EDFQD1 \input_weight_reg[5][64]  ( .D(data_in[64]), .E(n447), .CP(clk), .Q(
        \input_weight[5][64] ) );
  EDFQD1 \input_weight_reg[5][63]  ( .D(data_in[63]), .E(n447), .CP(clk), .Q(
        \input_weight[5][63] ) );
  EDFQD1 \input_weight_reg[5][62]  ( .D(data_in[62]), .E(n447), .CP(clk), .Q(
        \input_weight[5][62] ) );
  EDFQD1 \input_weight_reg[5][61]  ( .D(data_in[61]), .E(n447), .CP(clk), .Q(
        \input_weight[5][61] ) );
  EDFQD1 \input_weight_reg[5][60]  ( .D(data_in[60]), .E(n447), .CP(clk), .Q(
        \input_weight[5][60] ) );
  EDFQD1 \input_weight_reg[5][59]  ( .D(data_in[59]), .E(n447), .CP(clk), .Q(
        \input_weight[5][59] ) );
  EDFQD1 \input_weight_reg[5][58]  ( .D(data_in[58]), .E(n447), .CP(clk), .Q(
        \input_weight[5][58] ) );
  EDFQD1 \input_weight_reg[5][57]  ( .D(data_in[57]), .E(n447), .CP(clk), .Q(
        \input_weight[5][57] ) );
  EDFQD1 \input_weight_reg[5][56]  ( .D(data_in[56]), .E(n447), .CP(clk), .Q(
        \input_weight[5][56] ) );
  EDFQD1 \input_weight_reg[5][55]  ( .D(data_in[55]), .E(n447), .CP(clk), .Q(
        \input_weight[5][55] ) );
  EDFQD1 \input_weight_reg[5][54]  ( .D(data_in[54]), .E(n447), .CP(clk), .Q(
        \input_weight[5][54] ) );
  EDFQD1 \input_weight_reg[5][53]  ( .D(data_in[53]), .E(n447), .CP(clk), .Q(
        \input_weight[5][53] ) );
  EDFQD1 \input_weight_reg[5][52]  ( .D(data_in[52]), .E(n447), .CP(clk), .Q(
        \input_weight[5][52] ) );
  EDFQD1 \input_weight_reg[5][51]  ( .D(data_in[51]), .E(n446), .CP(clk), .Q(
        \input_weight[5][51] ) );
  EDFQD1 \input_weight_reg[5][50]  ( .D(data_in[50]), .E(n446), .CP(clk), .Q(
        \input_weight[5][50] ) );
  EDFQD1 \input_weight_reg[5][49]  ( .D(data_in[49]), .E(n446), .CP(clk), .Q(
        \input_weight[5][49] ) );
  EDFQD1 \input_weight_reg[5][48]  ( .D(data_in[48]), .E(n446), .CP(clk), .Q(
        \input_weight[5][48] ) );
  EDFQD1 \input_weight_reg[5][47]  ( .D(data_in[47]), .E(n446), .CP(clk), .Q(
        \input_weight[5][47] ) );
  EDFQD1 \input_weight_reg[5][46]  ( .D(data_in[46]), .E(n446), .CP(clk), .Q(
        \input_weight[5][46] ) );
  EDFQD1 \input_weight_reg[5][45]  ( .D(data_in[45]), .E(n446), .CP(clk), .Q(
        \input_weight[5][45] ) );
  EDFQD1 \input_weight_reg[5][44]  ( .D(data_in[44]), .E(n446), .CP(clk), .Q(
        \input_weight[5][44] ) );
  EDFQD1 \input_weight_reg[5][43]  ( .D(data_in[43]), .E(n446), .CP(clk), .Q(
        \input_weight[5][43] ) );
  EDFQD1 \input_weight_reg[5][42]  ( .D(data_in[42]), .E(n446), .CP(clk), .Q(
        \input_weight[5][42] ) );
  EDFQD1 \input_weight_reg[5][41]  ( .D(data_in[41]), .E(n446), .CP(clk), .Q(
        \input_weight[5][41] ) );
  EDFQD1 \input_weight_reg[5][40]  ( .D(data_in[40]), .E(n446), .CP(clk), .Q(
        \input_weight[5][40] ) );
  EDFQD1 \input_weight_reg[5][39]  ( .D(data_in[39]), .E(n446), .CP(clk), .Q(
        \input_weight[5][39] ) );
  EDFQD1 \input_weight_reg[5][38]  ( .D(data_in[38]), .E(n445), .CP(clk), .Q(
        \input_weight[5][38] ) );
  EDFQD1 \input_weight_reg[5][37]  ( .D(data_in[37]), .E(n445), .CP(clk), .Q(
        \input_weight[5][37] ) );
  EDFQD1 \input_weight_reg[5][36]  ( .D(data_in[36]), .E(n445), .CP(clk), .Q(
        \input_weight[5][36] ) );
  EDFQD1 \input_weight_reg[5][35]  ( .D(data_in[35]), .E(n445), .CP(clk), .Q(
        \input_weight[5][35] ) );
  EDFQD1 \input_weight_reg[5][34]  ( .D(data_in[34]), .E(n445), .CP(clk), .Q(
        \input_weight[5][34] ) );
  EDFQD1 \input_weight_reg[5][33]  ( .D(data_in[33]), .E(n445), .CP(clk), .Q(
        \input_weight[5][33] ) );
  EDFQD1 \input_weight_reg[5][32]  ( .D(data_in[32]), .E(n445), .CP(clk), .Q(
        \input_weight[5][32] ) );
  EDFQD1 \input_weight_reg[5][31]  ( .D(data_in[31]), .E(n445), .CP(clk), .Q(
        \input_weight[5][31] ) );
  EDFQD1 \input_weight_reg[5][30]  ( .D(data_in[30]), .E(n445), .CP(clk), .Q(
        \input_weight[5][30] ) );
  EDFQD1 \input_weight_reg[5][29]  ( .D(data_in[29]), .E(n445), .CP(clk), .Q(
        \input_weight[5][29] ) );
  EDFQD1 \input_weight_reg[5][28]  ( .D(data_in[28]), .E(n445), .CP(clk), .Q(
        \input_weight[5][28] ) );
  EDFQD1 \input_weight_reg[5][27]  ( .D(data_in[27]), .E(n445), .CP(clk), .Q(
        \input_weight[5][27] ) );
  EDFQD1 \input_weight_reg[5][26]  ( .D(data_in[26]), .E(n445), .CP(clk), .Q(
        \input_weight[5][26] ) );
  EDFQD1 \input_weight_reg[5][25]  ( .D(data_in[25]), .E(n444), .CP(clk), .Q(
        \input_weight[5][25] ) );
  EDFQD1 \input_weight_reg[5][24]  ( .D(data_in[24]), .E(n444), .CP(clk), .Q(
        \input_weight[5][24] ) );
  EDFQD1 \input_weight_reg[5][23]  ( .D(data_in[23]), .E(n444), .CP(clk), .Q(
        \input_weight[5][23] ) );
  EDFQD1 \input_weight_reg[5][22]  ( .D(data_in[22]), .E(n444), .CP(clk), .Q(
        \input_weight[5][22] ) );
  EDFQD1 \input_weight_reg[5][21]  ( .D(data_in[21]), .E(n444), .CP(clk), .Q(
        \input_weight[5][21] ) );
  EDFQD1 \input_weight_reg[5][20]  ( .D(data_in[20]), .E(n444), .CP(clk), .Q(
        \input_weight[5][20] ) );
  EDFQD1 \input_weight_reg[5][19]  ( .D(data_in[19]), .E(n444), .CP(clk), .Q(
        \input_weight[5][19] ) );
  EDFQD1 \input_weight_reg[5][18]  ( .D(data_in[18]), .E(n444), .CP(clk), .Q(
        \input_weight[5][18] ) );
  EDFQD1 \input_weight_reg[5][17]  ( .D(data_in[17]), .E(n444), .CP(clk), .Q(
        \input_weight[5][17] ) );
  EDFQD1 \input_weight_reg[5][16]  ( .D(data_in[16]), .E(n444), .CP(clk), .Q(
        \input_weight[5][16] ) );
  EDFQD1 \input_weight_reg[5][15]  ( .D(data_in[15]), .E(n444), .CP(clk), .Q(
        \input_weight[5][15] ) );
  EDFQD1 \input_weight_reg[5][14]  ( .D(data_in[14]), .E(n444), .CP(clk), .Q(
        \input_weight[5][14] ) );
  EDFQD1 \input_weight_reg[5][13]  ( .D(data_in[13]), .E(n444), .CP(clk), .Q(
        \input_weight[5][13] ) );
  EDFQD1 \input_weight_reg[5][12]  ( .D(data_in[12]), .E(n443), .CP(clk), .Q(
        \input_weight[5][12] ) );
  EDFQD1 \input_weight_reg[5][11]  ( .D(data_in[11]), .E(n443), .CP(clk), .Q(
        \input_weight[5][11] ) );
  EDFQD1 \input_weight_reg[5][10]  ( .D(data_in[10]), .E(n443), .CP(clk), .Q(
        \input_weight[5][10] ) );
  EDFQD1 \input_weight_reg[5][9]  ( .D(data_in[9]), .E(n443), .CP(clk), .Q(
        \input_weight[5][9] ) );
  EDFQD1 \input_weight_reg[5][8]  ( .D(data_in[8]), .E(n443), .CP(clk), .Q(
        \input_weight[5][8] ) );
  EDFQD1 \input_weight_reg[5][7]  ( .D(data_in[7]), .E(n443), .CP(clk), .Q(
        \input_weight[5][7] ) );
  EDFQD1 \input_weight_reg[5][6]  ( .D(data_in[6]), .E(n443), .CP(clk), .Q(
        \input_weight[5][6] ) );
  EDFQD1 \input_weight_reg[5][5]  ( .D(data_in[5]), .E(n443), .CP(clk), .Q(
        \input_weight[5][5] ) );
  EDFQD1 \input_weight_reg[5][4]  ( .D(data_in[4]), .E(n443), .CP(clk), .Q(
        \input_weight[5][4] ) );
  EDFQD1 \input_weight_reg[5][3]  ( .D(data_in[3]), .E(n443), .CP(clk), .Q(
        \input_weight[5][3] ) );
  EDFQD1 \input_weight_reg[5][2]  ( .D(data_in[2]), .E(n443), .CP(clk), .Q(
        \input_weight[5][2] ) );
  EDFQD1 \input_weight_reg[5][1]  ( .D(data_in[1]), .E(n443), .CP(clk), .Q(
        \input_weight[5][1] ) );
  EDFQD1 \input_weight_reg[5][0]  ( .D(data_in[0]), .E(n443), .CP(clk), .Q(
        \input_weight[5][0] ) );
  EDFQD1 \input_value_reg[1][99]  ( .D(data_in[99]), .E(n392), .CP(clk), .Q(
        \input_value[1][99] ) );
  EDFQD1 \input_value_reg[1][100]  ( .D(data_in[100]), .E(n392), .CP(clk), .Q(
        \input_value[1][100] ) );
  EDFQD1 \input_value_reg[1][101]  ( .D(data_in[101]), .E(n392), .CP(clk), .Q(
        \input_value[1][101] ) );
  EDFQD1 \input_value_reg[1][102]  ( .D(data_in[102]), .E(n392), .CP(clk), .Q(
        \input_value[1][102] ) );
  EDFQD1 \input_value_reg[1][103]  ( .D(data_in[103]), .E(n392), .CP(clk), .Q(
        \input_value[1][103] ) );
  EDFQD1 \input_value_reg[1][104]  ( .D(data_in[104]), .E(n392), .CP(clk), .Q(
        \input_value[1][104] ) );
  EDFQD1 \input_value_reg[1][105]  ( .D(data_in[105]), .E(n392), .CP(clk), .Q(
        \input_value[1][105] ) );
  EDFQD1 \input_value_reg[1][106]  ( .D(data_in[106]), .E(n392), .CP(clk), .Q(
        \input_value[1][106] ) );
  EDFQD1 \input_value_reg[1][107]  ( .D(data_in[107]), .E(n392), .CP(clk), .Q(
        \input_value[1][107] ) );
  EDFQD1 \input_value_reg[1][108]  ( .D(data_in[108]), .E(n392), .CP(clk), .Q(
        \input_value[1][108] ) );
  EDFQD1 \input_value_reg[1][109]  ( .D(data_in[109]), .E(n392), .CP(clk), .Q(
        \input_value[1][109] ) );
  EDFQD1 \input_value_reg[1][110]  ( .D(data_in[110]), .E(n391), .CP(clk), .Q(
        \input_value[1][110] ) );
  EDFQD1 \input_value_reg[1][111]  ( .D(data_in[111]), .E(n391), .CP(clk), .Q(
        \input_value[1][111] ) );
  EDFQD1 \input_value_reg[1][112]  ( .D(data_in[112]), .E(n391), .CP(clk), .Q(
        \input_value[1][112] ) );
  EDFQD1 \input_value_reg[1][113]  ( .D(data_in[113]), .E(n391), .CP(clk), .Q(
        \input_value[1][113] ) );
  EDFQD1 \input_value_reg[1][114]  ( .D(data_in[114]), .E(n391), .CP(clk), .Q(
        \input_value[1][114] ) );
  EDFQD1 \input_value_reg[1][115]  ( .D(data_in[115]), .E(n391), .CP(clk), .Q(
        \input_value[1][115] ) );
  EDFQD1 \input_value_reg[1][116]  ( .D(data_in[116]), .E(n391), .CP(clk), .Q(
        \input_value[1][116] ) );
  EDFQD1 \input_value_reg[1][117]  ( .D(data_in[117]), .E(n391), .CP(clk), .Q(
        \input_value[1][117] ) );
  EDFQD1 \input_value_reg[1][118]  ( .D(data_in[118]), .E(n391), .CP(clk), .Q(
        \input_value[1][118] ) );
  EDFQD1 \input_value_reg[1][119]  ( .D(data_in[119]), .E(n391), .CP(clk), .Q(
        \input_value[1][119] ) );
  EDFQD1 \input_value_reg[1][120]  ( .D(data_in[120]), .E(n391), .CP(clk), .Q(
        \input_value[1][120] ) );
  EDFQD1 \input_value_reg[1][121]  ( .D(data_in[121]), .E(n391), .CP(clk), .Q(
        \input_value[1][121] ) );
  EDFQD1 \input_value_reg[1][122]  ( .D(data_in[122]), .E(n391), .CP(clk), .Q(
        \input_value[1][122] ) );
  EDFQD1 \input_value_reg[1][123]  ( .D(data_in[123]), .E(n390), .CP(clk), .Q(
        \input_value[1][123] ) );
  EDFQD1 \input_value_reg[1][124]  ( .D(data_in[124]), .E(n390), .CP(clk), .Q(
        \input_value[1][124] ) );
  EDFQD1 \input_value_reg[1][125]  ( .D(data_in[125]), .E(n390), .CP(clk), .Q(
        \input_value[1][125] ) );
  EDFQD1 \input_value_reg[1][126]  ( .D(data_in[126]), .E(n390), .CP(clk), .Q(
        \input_value[1][126] ) );
  EDFQD1 \input_value_reg[1][127]  ( .D(data_in[127]), .E(n390), .CP(clk), .Q(
        \input_value[1][127] ) );
  EDFQD1 \input_value_reg[1][98]  ( .D(data_in[98]), .E(n390), .CP(clk), .Q(
        \input_value[1][98] ) );
  EDFQD1 \input_value_reg[1][97]  ( .D(data_in[97]), .E(n390), .CP(clk), .Q(
        \input_value[1][97] ) );
  EDFQD1 \input_value_reg[1][96]  ( .D(data_in[96]), .E(n390), .CP(clk), .Q(
        \input_value[1][96] ) );
  EDFQD1 \input_value_reg[1][95]  ( .D(data_in[95]), .E(n390), .CP(clk), .Q(
        \input_value[1][95] ) );
  EDFQD1 \input_value_reg[1][94]  ( .D(data_in[94]), .E(n390), .CP(clk), .Q(
        \input_value[1][94] ) );
  EDFQD1 \input_value_reg[1][93]  ( .D(data_in[93]), .E(n390), .CP(clk), .Q(
        \input_value[1][93] ) );
  EDFQD1 \input_value_reg[1][92]  ( .D(data_in[92]), .E(n390), .CP(clk), .Q(
        \input_value[1][92] ) );
  EDFQD1 \input_value_reg[1][91]  ( .D(data_in[91]), .E(n390), .CP(clk), .Q(
        \input_value[1][91] ) );
  EDFQD1 \input_value_reg[1][90]  ( .D(data_in[90]), .E(n389), .CP(clk), .Q(
        \input_value[1][90] ) );
  EDFQD1 \input_value_reg[1][89]  ( .D(data_in[89]), .E(n389), .CP(clk), .Q(
        \input_value[1][89] ) );
  EDFQD1 \input_value_reg[1][88]  ( .D(data_in[88]), .E(n389), .CP(clk), .Q(
        \input_value[1][88] ) );
  EDFQD1 \input_value_reg[1][87]  ( .D(data_in[87]), .E(n389), .CP(clk), .Q(
        \input_value[1][87] ) );
  EDFQD1 \input_value_reg[1][86]  ( .D(data_in[86]), .E(n389), .CP(clk), .Q(
        \input_value[1][86] ) );
  EDFQD1 \input_value_reg[1][85]  ( .D(data_in[85]), .E(n389), .CP(clk), .Q(
        \input_value[1][85] ) );
  EDFQD1 \input_value_reg[1][84]  ( .D(data_in[84]), .E(n389), .CP(clk), .Q(
        \input_value[1][84] ) );
  EDFQD1 \input_value_reg[1][83]  ( .D(data_in[83]), .E(n389), .CP(clk), .Q(
        \input_value[1][83] ) );
  EDFQD1 \input_value_reg[1][82]  ( .D(data_in[82]), .E(n389), .CP(clk), .Q(
        \input_value[1][82] ) );
  EDFQD1 \input_value_reg[1][81]  ( .D(data_in[81]), .E(n389), .CP(clk), .Q(
        \input_value[1][81] ) );
  EDFQD1 \input_value_reg[1][80]  ( .D(data_in[80]), .E(n389), .CP(clk), .Q(
        \input_value[1][80] ) );
  EDFQD1 \input_value_reg[1][79]  ( .D(data_in[79]), .E(n389), .CP(clk), .Q(
        \input_value[1][79] ) );
  EDFQD1 \input_value_reg[1][78]  ( .D(data_in[78]), .E(n389), .CP(clk), .Q(
        \input_value[1][78] ) );
  EDFQD1 \input_value_reg[1][77]  ( .D(data_in[77]), .E(n388), .CP(clk), .Q(
        \input_value[1][77] ) );
  EDFQD1 \input_value_reg[1][76]  ( .D(data_in[76]), .E(n388), .CP(clk), .Q(
        \input_value[1][76] ) );
  EDFQD1 \input_value_reg[1][75]  ( .D(data_in[75]), .E(n388), .CP(clk), .Q(
        \input_value[1][75] ) );
  EDFQD1 \input_value_reg[1][74]  ( .D(data_in[74]), .E(n388), .CP(clk), .Q(
        \input_value[1][74] ) );
  EDFQD1 \input_value_reg[1][73]  ( .D(data_in[73]), .E(n388), .CP(clk), .Q(
        \input_value[1][73] ) );
  EDFQD1 \input_value_reg[1][72]  ( .D(data_in[72]), .E(n388), .CP(clk), .Q(
        \input_value[1][72] ) );
  EDFQD1 \input_value_reg[1][71]  ( .D(data_in[71]), .E(n388), .CP(clk), .Q(
        \input_value[1][71] ) );
  EDFQD1 \input_value_reg[1][70]  ( .D(data_in[70]), .E(n388), .CP(clk), .Q(
        \input_value[1][70] ) );
  EDFQD1 \input_value_reg[1][69]  ( .D(data_in[69]), .E(n388), .CP(clk), .Q(
        \input_value[1][69] ) );
  EDFQD1 \input_value_reg[1][68]  ( .D(data_in[68]), .E(n388), .CP(clk), .Q(
        \input_value[1][68] ) );
  EDFQD1 \input_value_reg[1][67]  ( .D(data_in[67]), .E(n388), .CP(clk), .Q(
        \input_value[1][67] ) );
  EDFQD1 \input_value_reg[1][66]  ( .D(data_in[66]), .E(n388), .CP(clk), .Q(
        \input_value[1][66] ) );
  EDFQD1 \input_value_reg[1][65]  ( .D(data_in[65]), .E(n388), .CP(clk), .Q(
        \input_value[1][65] ) );
  EDFQD1 \input_value_reg[1][64]  ( .D(data_in[64]), .E(n387), .CP(clk), .Q(
        \input_value[1][64] ) );
  EDFQD1 \input_value_reg[1][63]  ( .D(data_in[63]), .E(n387), .CP(clk), .Q(
        \input_value[1][63] ) );
  EDFQD1 \input_value_reg[1][62]  ( .D(data_in[62]), .E(n387), .CP(clk), .Q(
        \input_value[1][62] ) );
  EDFQD1 \input_value_reg[1][61]  ( .D(data_in[61]), .E(n387), .CP(clk), .Q(
        \input_value[1][61] ) );
  EDFQD1 \input_value_reg[1][60]  ( .D(data_in[60]), .E(n387), .CP(clk), .Q(
        \input_value[1][60] ) );
  EDFQD1 \input_value_reg[1][59]  ( .D(data_in[59]), .E(n387), .CP(clk), .Q(
        \input_value[1][59] ) );
  EDFQD1 \input_value_reg[1][58]  ( .D(data_in[58]), .E(n387), .CP(clk), .Q(
        \input_value[1][58] ) );
  EDFQD1 \input_value_reg[1][57]  ( .D(data_in[57]), .E(n387), .CP(clk), .Q(
        \input_value[1][57] ) );
  EDFQD1 \input_value_reg[1][56]  ( .D(data_in[56]), .E(n387), .CP(clk), .Q(
        \input_value[1][56] ) );
  EDFQD1 \input_value_reg[1][55]  ( .D(data_in[55]), .E(n387), .CP(clk), .Q(
        \input_value[1][55] ) );
  EDFQD1 \input_value_reg[1][54]  ( .D(data_in[54]), .E(n387), .CP(clk), .Q(
        \input_value[1][54] ) );
  EDFQD1 \input_value_reg[1][53]  ( .D(data_in[53]), .E(n387), .CP(clk), .Q(
        \input_value[1][53] ) );
  EDFQD1 \input_value_reg[1][52]  ( .D(data_in[52]), .E(n387), .CP(clk), .Q(
        \input_value[1][52] ) );
  EDFQD1 \input_value_reg[1][51]  ( .D(data_in[51]), .E(n386), .CP(clk), .Q(
        \input_value[1][51] ) );
  EDFQD1 \input_value_reg[1][50]  ( .D(data_in[50]), .E(n386), .CP(clk), .Q(
        \input_value[1][50] ) );
  EDFQD1 \input_value_reg[1][49]  ( .D(data_in[49]), .E(n386), .CP(clk), .Q(
        \input_value[1][49] ) );
  EDFQD1 \input_value_reg[1][48]  ( .D(data_in[48]), .E(n386), .CP(clk), .Q(
        \input_value[1][48] ) );
  EDFQD1 \input_value_reg[1][47]  ( .D(data_in[47]), .E(n386), .CP(clk), .Q(
        \input_value[1][47] ) );
  EDFQD1 \input_value_reg[1][46]  ( .D(data_in[46]), .E(n386), .CP(clk), .Q(
        \input_value[1][46] ) );
  EDFQD1 \input_value_reg[1][45]  ( .D(data_in[45]), .E(n386), .CP(clk), .Q(
        \input_value[1][45] ) );
  EDFQD1 \input_value_reg[1][44]  ( .D(data_in[44]), .E(n386), .CP(clk), .Q(
        \input_value[1][44] ) );
  EDFQD1 \input_value_reg[1][43]  ( .D(data_in[43]), .E(n386), .CP(clk), .Q(
        \input_value[1][43] ) );
  EDFQD1 \input_value_reg[1][42]  ( .D(data_in[42]), .E(n386), .CP(clk), .Q(
        \input_value[1][42] ) );
  EDFQD1 \input_value_reg[1][41]  ( .D(data_in[41]), .E(n386), .CP(clk), .Q(
        \input_value[1][41] ) );
  EDFQD1 \input_value_reg[1][40]  ( .D(data_in[40]), .E(n386), .CP(clk), .Q(
        \input_value[1][40] ) );
  EDFQD1 \input_value_reg[1][39]  ( .D(data_in[39]), .E(n386), .CP(clk), .Q(
        \input_value[1][39] ) );
  EDFQD1 \input_value_reg[1][38]  ( .D(data_in[38]), .E(n385), .CP(clk), .Q(
        \input_value[1][38] ) );
  EDFQD1 \input_value_reg[1][37]  ( .D(data_in[37]), .E(n385), .CP(clk), .Q(
        \input_value[1][37] ) );
  EDFQD1 \input_value_reg[1][36]  ( .D(data_in[36]), .E(n385), .CP(clk), .Q(
        \input_value[1][36] ) );
  EDFQD1 \input_value_reg[1][35]  ( .D(data_in[35]), .E(n385), .CP(clk), .Q(
        \input_value[1][35] ) );
  EDFQD1 \input_value_reg[1][34]  ( .D(data_in[34]), .E(n385), .CP(clk), .Q(
        \input_value[1][34] ) );
  EDFQD1 \input_value_reg[1][33]  ( .D(data_in[33]), .E(n385), .CP(clk), .Q(
        \input_value[1][33] ) );
  EDFQD1 \input_value_reg[1][32]  ( .D(data_in[32]), .E(n385), .CP(clk), .Q(
        \input_value[1][32] ) );
  EDFQD1 \input_value_reg[1][31]  ( .D(data_in[31]), .E(n385), .CP(clk), .Q(
        \input_value[1][31] ) );
  EDFQD1 \input_value_reg[1][30]  ( .D(data_in[30]), .E(n385), .CP(clk), .Q(
        \input_value[1][30] ) );
  EDFQD1 \input_value_reg[1][29]  ( .D(data_in[29]), .E(n385), .CP(clk), .Q(
        \input_value[1][29] ) );
  EDFQD1 \input_value_reg[1][28]  ( .D(data_in[28]), .E(n385), .CP(clk), .Q(
        \input_value[1][28] ) );
  EDFQD1 \input_value_reg[1][27]  ( .D(data_in[27]), .E(n385), .CP(clk), .Q(
        \input_value[1][27] ) );
  EDFQD1 \input_value_reg[1][26]  ( .D(data_in[26]), .E(n385), .CP(clk), .Q(
        \input_value[1][26] ) );
  EDFQD1 \input_value_reg[1][25]  ( .D(data_in[25]), .E(n384), .CP(clk), .Q(
        \input_value[1][25] ) );
  EDFQD1 \input_value_reg[1][24]  ( .D(data_in[24]), .E(n384), .CP(clk), .Q(
        \input_value[1][24] ) );
  EDFQD1 \input_value_reg[1][23]  ( .D(data_in[23]), .E(n384), .CP(clk), .Q(
        \input_value[1][23] ) );
  EDFQD1 \input_value_reg[1][22]  ( .D(data_in[22]), .E(n384), .CP(clk), .Q(
        \input_value[1][22] ) );
  EDFQD1 \input_value_reg[1][21]  ( .D(data_in[21]), .E(n384), .CP(clk), .Q(
        \input_value[1][21] ) );
  EDFQD1 \input_value_reg[1][20]  ( .D(data_in[20]), .E(n384), .CP(clk), .Q(
        \input_value[1][20] ) );
  EDFQD1 \input_value_reg[1][19]  ( .D(data_in[19]), .E(n384), .CP(clk), .Q(
        \input_value[1][19] ) );
  EDFQD1 \input_value_reg[1][18]  ( .D(data_in[18]), .E(n384), .CP(clk), .Q(
        \input_value[1][18] ) );
  EDFQD1 \input_value_reg[1][17]  ( .D(data_in[17]), .E(n384), .CP(clk), .Q(
        \input_value[1][17] ) );
  EDFQD1 \input_value_reg[1][16]  ( .D(data_in[16]), .E(n384), .CP(clk), .Q(
        \input_value[1][16] ) );
  EDFQD1 \input_value_reg[1][15]  ( .D(data_in[15]), .E(n384), .CP(clk), .Q(
        \input_value[1][15] ) );
  EDFQD1 \input_value_reg[1][14]  ( .D(data_in[14]), .E(n384), .CP(clk), .Q(
        \input_value[1][14] ) );
  EDFQD1 \input_value_reg[1][13]  ( .D(data_in[13]), .E(n384), .CP(clk), .Q(
        \input_value[1][13] ) );
  EDFQD1 \input_value_reg[1][12]  ( .D(data_in[12]), .E(n383), .CP(clk), .Q(
        \input_value[1][12] ) );
  EDFQD1 \input_value_reg[1][11]  ( .D(data_in[11]), .E(n383), .CP(clk), .Q(
        \input_value[1][11] ) );
  EDFQD1 \input_value_reg[1][10]  ( .D(data_in[10]), .E(n383), .CP(clk), .Q(
        \input_value[1][10] ) );
  EDFQD1 \input_value_reg[1][9]  ( .D(data_in[9]), .E(n383), .CP(clk), .Q(
        \input_value[1][9] ) );
  EDFQD1 \input_value_reg[1][8]  ( .D(data_in[8]), .E(n383), .CP(clk), .Q(
        \input_value[1][8] ) );
  EDFQD1 \input_value_reg[1][7]  ( .D(data_in[7]), .E(n383), .CP(clk), .Q(
        \input_value[1][7] ) );
  EDFQD1 \input_value_reg[1][6]  ( .D(data_in[6]), .E(n383), .CP(clk), .Q(
        \input_value[1][6] ) );
  EDFQD1 \input_value_reg[1][5]  ( .D(data_in[5]), .E(n383), .CP(clk), .Q(
        \input_value[1][5] ) );
  EDFQD1 \input_value_reg[1][4]  ( .D(data_in[4]), .E(n383), .CP(clk), .Q(
        \input_value[1][4] ) );
  EDFQD1 \input_value_reg[1][3]  ( .D(data_in[3]), .E(n383), .CP(clk), .Q(
        \input_value[1][3] ) );
  EDFQD1 \input_value_reg[1][2]  ( .D(data_in[2]), .E(n383), .CP(clk), .Q(
        \input_value[1][2] ) );
  EDFQD1 \input_value_reg[1][1]  ( .D(data_in[1]), .E(n383), .CP(clk), .Q(
        \input_value[1][1] ) );
  EDFQD1 \input_value_reg[1][0]  ( .D(data_in[0]), .E(n383), .CP(clk), .Q(
        \input_value[1][0] ) );
  EDFQD1 \input_weight_reg[1][99]  ( .D(data_in[99]), .E(n512), .CP(clk), .Q(
        \input_weight[1][99] ) );
  EDFQD1 \input_weight_reg[1][100]  ( .D(data_in[100]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][100] ) );
  EDFQD1 \input_weight_reg[1][101]  ( .D(data_in[101]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][101] ) );
  EDFQD1 \input_weight_reg[1][102]  ( .D(data_in[102]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][102] ) );
  EDFQD1 \input_weight_reg[1][103]  ( .D(data_in[103]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][103] ) );
  EDFQD1 \input_weight_reg[1][104]  ( .D(data_in[104]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][104] ) );
  EDFQD1 \input_weight_reg[1][105]  ( .D(data_in[105]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][105] ) );
  EDFQD1 \input_weight_reg[1][106]  ( .D(data_in[106]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][106] ) );
  EDFQD1 \input_weight_reg[1][107]  ( .D(data_in[107]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][107] ) );
  EDFQD1 \input_weight_reg[1][108]  ( .D(data_in[108]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][108] ) );
  EDFQD1 \input_weight_reg[1][109]  ( .D(data_in[109]), .E(n512), .CP(clk), 
        .Q(\input_weight[1][109] ) );
  EDFQD1 \input_weight_reg[1][110]  ( .D(data_in[110]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][110] ) );
  EDFQD1 \input_weight_reg[1][111]  ( .D(data_in[111]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][111] ) );
  EDFQD1 \input_weight_reg[1][112]  ( .D(data_in[112]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][112] ) );
  EDFQD1 \input_weight_reg[1][113]  ( .D(data_in[113]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][113] ) );
  EDFQD1 \input_weight_reg[1][114]  ( .D(data_in[114]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][114] ) );
  EDFQD1 \input_weight_reg[1][115]  ( .D(data_in[115]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][115] ) );
  EDFQD1 \input_weight_reg[1][116]  ( .D(data_in[116]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][116] ) );
  EDFQD1 \input_weight_reg[1][117]  ( .D(data_in[117]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][117] ) );
  EDFQD1 \input_weight_reg[1][118]  ( .D(data_in[118]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][118] ) );
  EDFQD1 \input_weight_reg[1][119]  ( .D(data_in[119]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][119] ) );
  EDFQD1 \input_weight_reg[1][120]  ( .D(data_in[120]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][120] ) );
  EDFQD1 \input_weight_reg[1][121]  ( .D(data_in[121]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][121] ) );
  EDFQD1 \input_weight_reg[1][122]  ( .D(data_in[122]), .E(n511), .CP(clk), 
        .Q(\input_weight[1][122] ) );
  EDFQD1 \input_weight_reg[1][123]  ( .D(data_in[123]), .E(n510), .CP(clk), 
        .Q(\input_weight[1][123] ) );
  EDFQD1 \input_weight_reg[1][124]  ( .D(data_in[124]), .E(n510), .CP(clk), 
        .Q(\input_weight[1][124] ) );
  EDFQD1 \input_weight_reg[1][125]  ( .D(data_in[125]), .E(n510), .CP(clk), 
        .Q(\input_weight[1][125] ) );
  EDFQD1 \input_weight_reg[1][126]  ( .D(data_in[126]), .E(n510), .CP(clk), 
        .Q(\input_weight[1][126] ) );
  EDFQD1 \input_weight_reg[1][127]  ( .D(data_in[127]), .E(n510), .CP(clk), 
        .Q(\input_weight[1][127] ) );
  EDFQD1 \input_weight_reg[1][98]  ( .D(data_in[98]), .E(n510), .CP(clk), .Q(
        \input_weight[1][98] ) );
  EDFQD1 \input_weight_reg[1][97]  ( .D(data_in[97]), .E(n510), .CP(clk), .Q(
        \input_weight[1][97] ) );
  EDFQD1 \input_weight_reg[1][96]  ( .D(data_in[96]), .E(n510), .CP(clk), .Q(
        \input_weight[1][96] ) );
  EDFQD1 \input_weight_reg[1][95]  ( .D(data_in[95]), .E(n510), .CP(clk), .Q(
        \input_weight[1][95] ) );
  EDFQD1 \input_weight_reg[1][94]  ( .D(data_in[94]), .E(n510), .CP(clk), .Q(
        \input_weight[1][94] ) );
  EDFQD1 \input_weight_reg[1][93]  ( .D(data_in[93]), .E(n510), .CP(clk), .Q(
        \input_weight[1][93] ) );
  EDFQD1 \input_weight_reg[1][92]  ( .D(data_in[92]), .E(n510), .CP(clk), .Q(
        \input_weight[1][92] ) );
  EDFQD1 \input_weight_reg[1][91]  ( .D(data_in[91]), .E(n510), .CP(clk), .Q(
        \input_weight[1][91] ) );
  EDFQD1 \input_weight_reg[1][90]  ( .D(data_in[90]), .E(n509), .CP(clk), .Q(
        \input_weight[1][90] ) );
  EDFQD1 \input_weight_reg[1][89]  ( .D(data_in[89]), .E(n509), .CP(clk), .Q(
        \input_weight[1][89] ) );
  EDFQD1 \input_weight_reg[1][88]  ( .D(data_in[88]), .E(n509), .CP(clk), .Q(
        \input_weight[1][88] ) );
  EDFQD1 \input_weight_reg[1][87]  ( .D(data_in[87]), .E(n509), .CP(clk), .Q(
        \input_weight[1][87] ) );
  EDFQD1 \input_weight_reg[1][86]  ( .D(data_in[86]), .E(n509), .CP(clk), .Q(
        \input_weight[1][86] ) );
  EDFQD1 \input_weight_reg[1][85]  ( .D(data_in[85]), .E(n509), .CP(clk), .Q(
        \input_weight[1][85] ) );
  EDFQD1 \input_weight_reg[1][84]  ( .D(data_in[84]), .E(n509), .CP(clk), .Q(
        \input_weight[1][84] ) );
  EDFQD1 \input_weight_reg[1][83]  ( .D(data_in[83]), .E(n509), .CP(clk), .Q(
        \input_weight[1][83] ) );
  EDFQD1 \input_weight_reg[1][82]  ( .D(data_in[82]), .E(n509), .CP(clk), .Q(
        \input_weight[1][82] ) );
  EDFQD1 \input_weight_reg[1][81]  ( .D(data_in[81]), .E(n509), .CP(clk), .Q(
        \input_weight[1][81] ) );
  EDFQD1 \input_weight_reg[1][80]  ( .D(data_in[80]), .E(n509), .CP(clk), .Q(
        \input_weight[1][80] ) );
  EDFQD1 \input_weight_reg[1][79]  ( .D(data_in[79]), .E(n509), .CP(clk), .Q(
        \input_weight[1][79] ) );
  EDFQD1 \input_weight_reg[1][78]  ( .D(data_in[78]), .E(n509), .CP(clk), .Q(
        \input_weight[1][78] ) );
  EDFQD1 \input_weight_reg[1][77]  ( .D(data_in[77]), .E(n508), .CP(clk), .Q(
        \input_weight[1][77] ) );
  EDFQD1 \input_weight_reg[1][76]  ( .D(data_in[76]), .E(n508), .CP(clk), .Q(
        \input_weight[1][76] ) );
  EDFQD1 \input_weight_reg[1][75]  ( .D(data_in[75]), .E(n508), .CP(clk), .Q(
        \input_weight[1][75] ) );
  EDFQD1 \input_weight_reg[1][74]  ( .D(data_in[74]), .E(n508), .CP(clk), .Q(
        \input_weight[1][74] ) );
  EDFQD1 \input_weight_reg[1][73]  ( .D(data_in[73]), .E(n508), .CP(clk), .Q(
        \input_weight[1][73] ) );
  EDFQD1 \input_weight_reg[1][72]  ( .D(data_in[72]), .E(n508), .CP(clk), .Q(
        \input_weight[1][72] ) );
  EDFQD1 \input_weight_reg[1][71]  ( .D(data_in[71]), .E(n508), .CP(clk), .Q(
        \input_weight[1][71] ) );
  EDFQD1 \input_weight_reg[1][70]  ( .D(data_in[70]), .E(n508), .CP(clk), .Q(
        \input_weight[1][70] ) );
  EDFQD1 \input_weight_reg[1][69]  ( .D(data_in[69]), .E(n508), .CP(clk), .Q(
        \input_weight[1][69] ) );
  EDFQD1 \input_weight_reg[1][68]  ( .D(data_in[68]), .E(n508), .CP(clk), .Q(
        \input_weight[1][68] ) );
  EDFQD1 \input_weight_reg[1][67]  ( .D(data_in[67]), .E(n508), .CP(clk), .Q(
        \input_weight[1][67] ) );
  EDFQD1 \input_weight_reg[1][66]  ( .D(data_in[66]), .E(n508), .CP(clk), .Q(
        \input_weight[1][66] ) );
  EDFQD1 \input_weight_reg[1][65]  ( .D(data_in[65]), .E(n508), .CP(clk), .Q(
        \input_weight[1][65] ) );
  EDFQD1 \input_weight_reg[1][64]  ( .D(data_in[64]), .E(n507), .CP(clk), .Q(
        \input_weight[1][64] ) );
  EDFQD1 \input_weight_reg[1][63]  ( .D(data_in[63]), .E(n507), .CP(clk), .Q(
        \input_weight[1][63] ) );
  EDFQD1 \input_weight_reg[1][62]  ( .D(data_in[62]), .E(n507), .CP(clk), .Q(
        \input_weight[1][62] ) );
  EDFQD1 \input_weight_reg[1][61]  ( .D(data_in[61]), .E(n507), .CP(clk), .Q(
        \input_weight[1][61] ) );
  EDFQD1 \input_weight_reg[1][60]  ( .D(data_in[60]), .E(n507), .CP(clk), .Q(
        \input_weight[1][60] ) );
  EDFQD1 \input_weight_reg[1][59]  ( .D(data_in[59]), .E(n507), .CP(clk), .Q(
        \input_weight[1][59] ) );
  EDFQD1 \input_weight_reg[1][58]  ( .D(data_in[58]), .E(n507), .CP(clk), .Q(
        \input_weight[1][58] ) );
  EDFQD1 \input_weight_reg[1][57]  ( .D(data_in[57]), .E(n507), .CP(clk), .Q(
        \input_weight[1][57] ) );
  EDFQD1 \input_weight_reg[1][56]  ( .D(data_in[56]), .E(n507), .CP(clk), .Q(
        \input_weight[1][56] ) );
  EDFQD1 \input_weight_reg[1][55]  ( .D(data_in[55]), .E(n507), .CP(clk), .Q(
        \input_weight[1][55] ) );
  EDFQD1 \input_weight_reg[1][54]  ( .D(data_in[54]), .E(n507), .CP(clk), .Q(
        \input_weight[1][54] ) );
  EDFQD1 \input_weight_reg[1][53]  ( .D(data_in[53]), .E(n507), .CP(clk), .Q(
        \input_weight[1][53] ) );
  EDFQD1 \input_weight_reg[1][52]  ( .D(data_in[52]), .E(n507), .CP(clk), .Q(
        \input_weight[1][52] ) );
  EDFQD1 \input_weight_reg[1][51]  ( .D(data_in[51]), .E(n506), .CP(clk), .Q(
        \input_weight[1][51] ) );
  EDFQD1 \input_weight_reg[1][50]  ( .D(data_in[50]), .E(n506), .CP(clk), .Q(
        \input_weight[1][50] ) );
  EDFQD1 \input_weight_reg[1][49]  ( .D(data_in[49]), .E(n506), .CP(clk), .Q(
        \input_weight[1][49] ) );
  EDFQD1 \input_weight_reg[1][48]  ( .D(data_in[48]), .E(n506), .CP(clk), .Q(
        \input_weight[1][48] ) );
  EDFQD1 \input_weight_reg[1][47]  ( .D(data_in[47]), .E(n506), .CP(clk), .Q(
        \input_weight[1][47] ) );
  EDFQD1 \input_weight_reg[1][46]  ( .D(data_in[46]), .E(n506), .CP(clk), .Q(
        \input_weight[1][46] ) );
  EDFQD1 \input_weight_reg[1][45]  ( .D(data_in[45]), .E(n506), .CP(clk), .Q(
        \input_weight[1][45] ) );
  EDFQD1 \input_weight_reg[1][44]  ( .D(data_in[44]), .E(n506), .CP(clk), .Q(
        \input_weight[1][44] ) );
  EDFQD1 \input_weight_reg[1][43]  ( .D(data_in[43]), .E(n506), .CP(clk), .Q(
        \input_weight[1][43] ) );
  EDFQD1 \input_weight_reg[1][42]  ( .D(data_in[42]), .E(n506), .CP(clk), .Q(
        \input_weight[1][42] ) );
  EDFQD1 \input_weight_reg[1][41]  ( .D(data_in[41]), .E(n506), .CP(clk), .Q(
        \input_weight[1][41] ) );
  EDFQD1 \input_weight_reg[1][40]  ( .D(data_in[40]), .E(n506), .CP(clk), .Q(
        \input_weight[1][40] ) );
  EDFQD1 \input_weight_reg[1][39]  ( .D(data_in[39]), .E(n506), .CP(clk), .Q(
        \input_weight[1][39] ) );
  EDFQD1 \input_weight_reg[1][38]  ( .D(data_in[38]), .E(n505), .CP(clk), .Q(
        \input_weight[1][38] ) );
  EDFQD1 \input_weight_reg[1][37]  ( .D(data_in[37]), .E(n505), .CP(clk), .Q(
        \input_weight[1][37] ) );
  EDFQD1 \input_weight_reg[1][36]  ( .D(data_in[36]), .E(n505), .CP(clk), .Q(
        \input_weight[1][36] ) );
  EDFQD1 \input_weight_reg[1][35]  ( .D(data_in[35]), .E(n505), .CP(clk), .Q(
        \input_weight[1][35] ) );
  EDFQD1 \input_weight_reg[1][34]  ( .D(data_in[34]), .E(n505), .CP(clk), .Q(
        \input_weight[1][34] ) );
  EDFQD1 \input_weight_reg[1][33]  ( .D(data_in[33]), .E(n505), .CP(clk), .Q(
        \input_weight[1][33] ) );
  EDFQD1 \input_weight_reg[1][32]  ( .D(data_in[32]), .E(n505), .CP(clk), .Q(
        \input_weight[1][32] ) );
  EDFQD1 \input_weight_reg[1][31]  ( .D(data_in[31]), .E(n505), .CP(clk), .Q(
        \input_weight[1][31] ) );
  EDFQD1 \input_weight_reg[1][30]  ( .D(data_in[30]), .E(n505), .CP(clk), .Q(
        \input_weight[1][30] ) );
  EDFQD1 \input_weight_reg[1][29]  ( .D(data_in[29]), .E(n505), .CP(clk), .Q(
        \input_weight[1][29] ) );
  EDFQD1 \input_weight_reg[1][28]  ( .D(data_in[28]), .E(n505), .CP(clk), .Q(
        \input_weight[1][28] ) );
  EDFQD1 \input_weight_reg[1][27]  ( .D(data_in[27]), .E(n505), .CP(clk), .Q(
        \input_weight[1][27] ) );
  EDFQD1 \input_weight_reg[1][26]  ( .D(data_in[26]), .E(n505), .CP(clk), .Q(
        \input_weight[1][26] ) );
  EDFQD1 \input_weight_reg[1][25]  ( .D(data_in[25]), .E(n504), .CP(clk), .Q(
        \input_weight[1][25] ) );
  EDFQD1 \input_weight_reg[1][24]  ( .D(data_in[24]), .E(n504), .CP(clk), .Q(
        \input_weight[1][24] ) );
  EDFQD1 \input_weight_reg[1][23]  ( .D(data_in[23]), .E(n504), .CP(clk), .Q(
        \input_weight[1][23] ) );
  EDFQD1 \input_weight_reg[1][22]  ( .D(data_in[22]), .E(n504), .CP(clk), .Q(
        \input_weight[1][22] ) );
  EDFQD1 \input_weight_reg[1][21]  ( .D(data_in[21]), .E(n504), .CP(clk), .Q(
        \input_weight[1][21] ) );
  EDFQD1 \input_weight_reg[1][20]  ( .D(data_in[20]), .E(n504), .CP(clk), .Q(
        \input_weight[1][20] ) );
  EDFQD1 \input_weight_reg[1][19]  ( .D(data_in[19]), .E(n504), .CP(clk), .Q(
        \input_weight[1][19] ) );
  EDFQD1 \input_weight_reg[1][18]  ( .D(data_in[18]), .E(n504), .CP(clk), .Q(
        \input_weight[1][18] ) );
  EDFQD1 \input_weight_reg[1][17]  ( .D(data_in[17]), .E(n504), .CP(clk), .Q(
        \input_weight[1][17] ) );
  EDFQD1 \input_weight_reg[1][16]  ( .D(data_in[16]), .E(n504), .CP(clk), .Q(
        \input_weight[1][16] ) );
  EDFQD1 \input_weight_reg[1][15]  ( .D(data_in[15]), .E(n504), .CP(clk), .Q(
        \input_weight[1][15] ) );
  EDFQD1 \input_weight_reg[1][14]  ( .D(data_in[14]), .E(n504), .CP(clk), .Q(
        \input_weight[1][14] ) );
  EDFQD1 \input_weight_reg[1][13]  ( .D(data_in[13]), .E(n504), .CP(clk), .Q(
        \input_weight[1][13] ) );
  EDFQD1 \input_weight_reg[1][12]  ( .D(data_in[12]), .E(n503), .CP(clk), .Q(
        \input_weight[1][12] ) );
  EDFQD1 \input_weight_reg[1][11]  ( .D(data_in[11]), .E(n503), .CP(clk), .Q(
        \input_weight[1][11] ) );
  EDFQD1 \input_weight_reg[1][10]  ( .D(data_in[10]), .E(n503), .CP(clk), .Q(
        \input_weight[1][10] ) );
  EDFQD1 \input_weight_reg[1][9]  ( .D(data_in[9]), .E(n503), .CP(clk), .Q(
        \input_weight[1][9] ) );
  EDFQD1 \input_weight_reg[1][8]  ( .D(data_in[8]), .E(n503), .CP(clk), .Q(
        \input_weight[1][8] ) );
  EDFQD1 \input_weight_reg[1][7]  ( .D(data_in[7]), .E(n503), .CP(clk), .Q(
        \input_weight[1][7] ) );
  EDFQD1 \input_weight_reg[1][6]  ( .D(data_in[6]), .E(n503), .CP(clk), .Q(
        \input_weight[1][6] ) );
  EDFQD1 \input_weight_reg[1][5]  ( .D(data_in[5]), .E(n503), .CP(clk), .Q(
        \input_weight[1][5] ) );
  EDFQD1 \input_weight_reg[1][4]  ( .D(data_in[4]), .E(n503), .CP(clk), .Q(
        \input_weight[1][4] ) );
  EDFQD1 \input_weight_reg[1][3]  ( .D(data_in[3]), .E(n503), .CP(clk), .Q(
        \input_weight[1][3] ) );
  EDFQD1 \input_weight_reg[1][2]  ( .D(data_in[2]), .E(n503), .CP(clk), .Q(
        \input_weight[1][2] ) );
  EDFQD1 \input_weight_reg[1][1]  ( .D(data_in[1]), .E(n503), .CP(clk), .Q(
        \input_weight[1][1] ) );
  EDFQD1 \input_weight_reg[1][0]  ( .D(data_in[0]), .E(n503), .CP(clk), .Q(
        \input_weight[1][0] ) );
  EDFQD1 \input_value_reg[3][99]  ( .D(data_in[99]), .E(n362), .CP(clk), .Q(
        \input_value[3][99] ) );
  EDFQD1 \input_value_reg[3][100]  ( .D(data_in[100]), .E(n362), .CP(clk), .Q(
        \input_value[3][100] ) );
  EDFQD1 \input_value_reg[3][101]  ( .D(data_in[101]), .E(n362), .CP(clk), .Q(
        \input_value[3][101] ) );
  EDFQD1 \input_value_reg[3][102]  ( .D(data_in[102]), .E(n362), .CP(clk), .Q(
        \input_value[3][102] ) );
  EDFQD1 \input_value_reg[3][103]  ( .D(data_in[103]), .E(n362), .CP(clk), .Q(
        \input_value[3][103] ) );
  EDFQD1 \input_value_reg[3][104]  ( .D(data_in[104]), .E(n362), .CP(clk), .Q(
        \input_value[3][104] ) );
  EDFQD1 \input_value_reg[3][105]  ( .D(data_in[105]), .E(n362), .CP(clk), .Q(
        \input_value[3][105] ) );
  EDFQD1 \input_value_reg[3][106]  ( .D(data_in[106]), .E(n362), .CP(clk), .Q(
        \input_value[3][106] ) );
  EDFQD1 \input_value_reg[3][107]  ( .D(data_in[107]), .E(n362), .CP(clk), .Q(
        \input_value[3][107] ) );
  EDFQD1 \input_value_reg[3][108]  ( .D(data_in[108]), .E(n362), .CP(clk), .Q(
        \input_value[3][108] ) );
  EDFQD1 \input_value_reg[3][109]  ( .D(data_in[109]), .E(n362), .CP(clk), .Q(
        \input_value[3][109] ) );
  EDFQD1 \input_value_reg[3][110]  ( .D(data_in[110]), .E(n361), .CP(clk), .Q(
        \input_value[3][110] ) );
  EDFQD1 \input_value_reg[3][111]  ( .D(data_in[111]), .E(n361), .CP(clk), .Q(
        \input_value[3][111] ) );
  EDFQD1 \input_value_reg[3][112]  ( .D(data_in[112]), .E(n361), .CP(clk), .Q(
        \input_value[3][112] ) );
  EDFQD1 \input_value_reg[3][113]  ( .D(data_in[113]), .E(n361), .CP(clk), .Q(
        \input_value[3][113] ) );
  EDFQD1 \input_value_reg[3][114]  ( .D(data_in[114]), .E(n361), .CP(clk), .Q(
        \input_value[3][114] ) );
  EDFQD1 \input_value_reg[3][115]  ( .D(data_in[115]), .E(n361), .CP(clk), .Q(
        \input_value[3][115] ) );
  EDFQD1 \input_value_reg[3][116]  ( .D(data_in[116]), .E(n361), .CP(clk), .Q(
        \input_value[3][116] ) );
  EDFQD1 \input_value_reg[3][117]  ( .D(data_in[117]), .E(n361), .CP(clk), .Q(
        \input_value[3][117] ) );
  EDFQD1 \input_value_reg[3][118]  ( .D(data_in[118]), .E(n361), .CP(clk), .Q(
        \input_value[3][118] ) );
  EDFQD1 \input_value_reg[3][119]  ( .D(data_in[119]), .E(n361), .CP(clk), .Q(
        \input_value[3][119] ) );
  EDFQD1 \input_value_reg[3][120]  ( .D(data_in[120]), .E(n361), .CP(clk), .Q(
        \input_value[3][120] ) );
  EDFQD1 \input_value_reg[3][121]  ( .D(data_in[121]), .E(n361), .CP(clk), .Q(
        \input_value[3][121] ) );
  EDFQD1 \input_value_reg[3][122]  ( .D(data_in[122]), .E(n361), .CP(clk), .Q(
        \input_value[3][122] ) );
  EDFQD1 \input_value_reg[3][123]  ( .D(data_in[123]), .E(n360), .CP(clk), .Q(
        \input_value[3][123] ) );
  EDFQD1 \input_value_reg[3][124]  ( .D(data_in[124]), .E(n360), .CP(clk), .Q(
        \input_value[3][124] ) );
  EDFQD1 \input_value_reg[3][125]  ( .D(data_in[125]), .E(n360), .CP(clk), .Q(
        \input_value[3][125] ) );
  EDFQD1 \input_value_reg[3][126]  ( .D(data_in[126]), .E(n360), .CP(clk), .Q(
        \input_value[3][126] ) );
  EDFQD1 \input_value_reg[3][127]  ( .D(data_in[127]), .E(n360), .CP(clk), .Q(
        \input_value[3][127] ) );
  EDFQD1 \input_value_reg[3][98]  ( .D(data_in[98]), .E(n360), .CP(clk), .Q(
        \input_value[3][98] ) );
  EDFQD1 \input_value_reg[3][97]  ( .D(data_in[97]), .E(n360), .CP(clk), .Q(
        \input_value[3][97] ) );
  EDFQD1 \input_value_reg[3][96]  ( .D(data_in[96]), .E(n360), .CP(clk), .Q(
        \input_value[3][96] ) );
  EDFQD1 \input_value_reg[3][95]  ( .D(data_in[95]), .E(n360), .CP(clk), .Q(
        \input_value[3][95] ) );
  EDFQD1 \input_value_reg[3][94]  ( .D(data_in[94]), .E(n360), .CP(clk), .Q(
        \input_value[3][94] ) );
  EDFQD1 \input_value_reg[3][93]  ( .D(data_in[93]), .E(n360), .CP(clk), .Q(
        \input_value[3][93] ) );
  EDFQD1 \input_value_reg[3][92]  ( .D(data_in[92]), .E(n360), .CP(clk), .Q(
        \input_value[3][92] ) );
  EDFQD1 \input_value_reg[3][91]  ( .D(data_in[91]), .E(n360), .CP(clk), .Q(
        \input_value[3][91] ) );
  EDFQD1 \input_value_reg[3][90]  ( .D(data_in[90]), .E(n359), .CP(clk), .Q(
        \input_value[3][90] ) );
  EDFQD1 \input_value_reg[3][89]  ( .D(data_in[89]), .E(n359), .CP(clk), .Q(
        \input_value[3][89] ) );
  EDFQD1 \input_value_reg[3][88]  ( .D(data_in[88]), .E(n359), .CP(clk), .Q(
        \input_value[3][88] ) );
  EDFQD1 \input_value_reg[3][87]  ( .D(data_in[87]), .E(n359), .CP(clk), .Q(
        \input_value[3][87] ) );
  EDFQD1 \input_value_reg[3][86]  ( .D(data_in[86]), .E(n359), .CP(clk), .Q(
        \input_value[3][86] ) );
  EDFQD1 \input_value_reg[3][85]  ( .D(data_in[85]), .E(n359), .CP(clk), .Q(
        \input_value[3][85] ) );
  EDFQD1 \input_value_reg[3][84]  ( .D(data_in[84]), .E(n359), .CP(clk), .Q(
        \input_value[3][84] ) );
  EDFQD1 \input_value_reg[3][83]  ( .D(data_in[83]), .E(n359), .CP(clk), .Q(
        \input_value[3][83] ) );
  EDFQD1 \input_value_reg[3][82]  ( .D(data_in[82]), .E(n359), .CP(clk), .Q(
        \input_value[3][82] ) );
  EDFQD1 \input_value_reg[3][81]  ( .D(data_in[81]), .E(n359), .CP(clk), .Q(
        \input_value[3][81] ) );
  EDFQD1 \input_value_reg[3][80]  ( .D(data_in[80]), .E(n359), .CP(clk), .Q(
        \input_value[3][80] ) );
  EDFQD1 \input_value_reg[3][79]  ( .D(data_in[79]), .E(n359), .CP(clk), .Q(
        \input_value[3][79] ) );
  EDFQD1 \input_value_reg[3][78]  ( .D(data_in[78]), .E(n359), .CP(clk), .Q(
        \input_value[3][78] ) );
  EDFQD1 \input_value_reg[3][77]  ( .D(data_in[77]), .E(n358), .CP(clk), .Q(
        \input_value[3][77] ) );
  EDFQD1 \input_value_reg[3][76]  ( .D(data_in[76]), .E(n358), .CP(clk), .Q(
        \input_value[3][76] ) );
  EDFQD1 \input_value_reg[3][75]  ( .D(data_in[75]), .E(n358), .CP(clk), .Q(
        \input_value[3][75] ) );
  EDFQD1 \input_value_reg[3][74]  ( .D(data_in[74]), .E(n358), .CP(clk), .Q(
        \input_value[3][74] ) );
  EDFQD1 \input_value_reg[3][73]  ( .D(data_in[73]), .E(n358), .CP(clk), .Q(
        \input_value[3][73] ) );
  EDFQD1 \input_value_reg[3][72]  ( .D(data_in[72]), .E(n358), .CP(clk), .Q(
        \input_value[3][72] ) );
  EDFQD1 \input_value_reg[3][71]  ( .D(data_in[71]), .E(n358), .CP(clk), .Q(
        \input_value[3][71] ) );
  EDFQD1 \input_value_reg[3][70]  ( .D(data_in[70]), .E(n358), .CP(clk), .Q(
        \input_value[3][70] ) );
  EDFQD1 \input_value_reg[3][69]  ( .D(data_in[69]), .E(n358), .CP(clk), .Q(
        \input_value[3][69] ) );
  EDFQD1 \input_value_reg[3][68]  ( .D(data_in[68]), .E(n358), .CP(clk), .Q(
        \input_value[3][68] ) );
  EDFQD1 \input_value_reg[3][67]  ( .D(data_in[67]), .E(n358), .CP(clk), .Q(
        \input_value[3][67] ) );
  EDFQD1 \input_value_reg[3][66]  ( .D(data_in[66]), .E(n358), .CP(clk), .Q(
        \input_value[3][66] ) );
  EDFQD1 \input_value_reg[3][65]  ( .D(data_in[65]), .E(n358), .CP(clk), .Q(
        \input_value[3][65] ) );
  EDFQD1 \input_value_reg[3][64]  ( .D(data_in[64]), .E(n357), .CP(clk), .Q(
        \input_value[3][64] ) );
  EDFQD1 \input_value_reg[3][63]  ( .D(data_in[63]), .E(n357), .CP(clk), .Q(
        \input_value[3][63] ) );
  EDFQD1 \input_value_reg[3][62]  ( .D(data_in[62]), .E(n357), .CP(clk), .Q(
        \input_value[3][62] ) );
  EDFQD1 \input_value_reg[3][61]  ( .D(data_in[61]), .E(n357), .CP(clk), .Q(
        \input_value[3][61] ) );
  EDFQD1 \input_value_reg[3][60]  ( .D(data_in[60]), .E(n357), .CP(clk), .Q(
        \input_value[3][60] ) );
  EDFQD1 \input_value_reg[3][59]  ( .D(data_in[59]), .E(n357), .CP(clk), .Q(
        \input_value[3][59] ) );
  EDFQD1 \input_value_reg[3][58]  ( .D(data_in[58]), .E(n357), .CP(clk), .Q(
        \input_value[3][58] ) );
  EDFQD1 \input_value_reg[3][57]  ( .D(data_in[57]), .E(n357), .CP(clk), .Q(
        \input_value[3][57] ) );
  EDFQD1 \input_value_reg[3][56]  ( .D(data_in[56]), .E(n357), .CP(clk), .Q(
        \input_value[3][56] ) );
  EDFQD1 \input_value_reg[3][55]  ( .D(data_in[55]), .E(n357), .CP(clk), .Q(
        \input_value[3][55] ) );
  EDFQD1 \input_value_reg[3][54]  ( .D(data_in[54]), .E(n357), .CP(clk), .Q(
        \input_value[3][54] ) );
  EDFQD1 \input_value_reg[3][53]  ( .D(data_in[53]), .E(n357), .CP(clk), .Q(
        \input_value[3][53] ) );
  EDFQD1 \input_value_reg[3][52]  ( .D(data_in[52]), .E(n357), .CP(clk), .Q(
        \input_value[3][52] ) );
  EDFQD1 \input_value_reg[3][51]  ( .D(data_in[51]), .E(n356), .CP(clk), .Q(
        \input_value[3][51] ) );
  EDFQD1 \input_value_reg[3][50]  ( .D(data_in[50]), .E(n356), .CP(clk), .Q(
        \input_value[3][50] ) );
  EDFQD1 \input_value_reg[3][49]  ( .D(data_in[49]), .E(n356), .CP(clk), .Q(
        \input_value[3][49] ) );
  EDFQD1 \input_value_reg[3][48]  ( .D(data_in[48]), .E(n356), .CP(clk), .Q(
        \input_value[3][48] ) );
  EDFQD1 \input_value_reg[3][47]  ( .D(data_in[47]), .E(n356), .CP(clk), .Q(
        \input_value[3][47] ) );
  EDFQD1 \input_value_reg[3][46]  ( .D(data_in[46]), .E(n356), .CP(clk), .Q(
        \input_value[3][46] ) );
  EDFQD1 \input_value_reg[3][45]  ( .D(data_in[45]), .E(n356), .CP(clk), .Q(
        \input_value[3][45] ) );
  EDFQD1 \input_value_reg[3][44]  ( .D(data_in[44]), .E(n356), .CP(clk), .Q(
        \input_value[3][44] ) );
  EDFQD1 \input_value_reg[3][43]  ( .D(data_in[43]), .E(n356), .CP(clk), .Q(
        \input_value[3][43] ) );
  EDFQD1 \input_value_reg[3][42]  ( .D(data_in[42]), .E(n356), .CP(clk), .Q(
        \input_value[3][42] ) );
  EDFQD1 \input_value_reg[3][41]  ( .D(data_in[41]), .E(n356), .CP(clk), .Q(
        \input_value[3][41] ) );
  EDFQD1 \input_value_reg[3][40]  ( .D(data_in[40]), .E(n356), .CP(clk), .Q(
        \input_value[3][40] ) );
  EDFQD1 \input_value_reg[3][39]  ( .D(data_in[39]), .E(n356), .CP(clk), .Q(
        \input_value[3][39] ) );
  EDFQD1 \input_value_reg[3][38]  ( .D(data_in[38]), .E(n355), .CP(clk), .Q(
        \input_value[3][38] ) );
  EDFQD1 \input_value_reg[3][37]  ( .D(data_in[37]), .E(n355), .CP(clk), .Q(
        \input_value[3][37] ) );
  EDFQD1 \input_value_reg[3][36]  ( .D(data_in[36]), .E(n355), .CP(clk), .Q(
        \input_value[3][36] ) );
  EDFQD1 \input_value_reg[3][35]  ( .D(data_in[35]), .E(n355), .CP(clk), .Q(
        \input_value[3][35] ) );
  EDFQD1 \input_value_reg[3][34]  ( .D(data_in[34]), .E(n355), .CP(clk), .Q(
        \input_value[3][34] ) );
  EDFQD1 \input_value_reg[3][33]  ( .D(data_in[33]), .E(n355), .CP(clk), .Q(
        \input_value[3][33] ) );
  EDFQD1 \input_value_reg[3][32]  ( .D(data_in[32]), .E(n355), .CP(clk), .Q(
        \input_value[3][32] ) );
  EDFQD1 \input_value_reg[3][31]  ( .D(data_in[31]), .E(n355), .CP(clk), .Q(
        \input_value[3][31] ) );
  EDFQD1 \input_value_reg[3][30]  ( .D(data_in[30]), .E(n355), .CP(clk), .Q(
        \input_value[3][30] ) );
  EDFQD1 \input_value_reg[3][29]  ( .D(data_in[29]), .E(n355), .CP(clk), .Q(
        \input_value[3][29] ) );
  EDFQD1 \input_value_reg[3][28]  ( .D(data_in[28]), .E(n355), .CP(clk), .Q(
        \input_value[3][28] ) );
  EDFQD1 \input_value_reg[3][27]  ( .D(data_in[27]), .E(n355), .CP(clk), .Q(
        \input_value[3][27] ) );
  EDFQD1 \input_value_reg[3][26]  ( .D(data_in[26]), .E(n355), .CP(clk), .Q(
        \input_value[3][26] ) );
  EDFQD1 \input_value_reg[3][25]  ( .D(data_in[25]), .E(n354), .CP(clk), .Q(
        \input_value[3][25] ) );
  EDFQD1 \input_value_reg[3][24]  ( .D(data_in[24]), .E(n354), .CP(clk), .Q(
        \input_value[3][24] ) );
  EDFQD1 \input_value_reg[3][23]  ( .D(data_in[23]), .E(n354), .CP(clk), .Q(
        \input_value[3][23] ) );
  EDFQD1 \input_value_reg[3][22]  ( .D(data_in[22]), .E(n354), .CP(clk), .Q(
        \input_value[3][22] ) );
  EDFQD1 \input_value_reg[3][21]  ( .D(data_in[21]), .E(n354), .CP(clk), .Q(
        \input_value[3][21] ) );
  EDFQD1 \input_value_reg[3][20]  ( .D(data_in[20]), .E(n354), .CP(clk), .Q(
        \input_value[3][20] ) );
  EDFQD1 \input_value_reg[3][19]  ( .D(data_in[19]), .E(n354), .CP(clk), .Q(
        \input_value[3][19] ) );
  EDFQD1 \input_value_reg[3][18]  ( .D(data_in[18]), .E(n354), .CP(clk), .Q(
        \input_value[3][18] ) );
  EDFQD1 \input_value_reg[3][17]  ( .D(data_in[17]), .E(n354), .CP(clk), .Q(
        \input_value[3][17] ) );
  EDFQD1 \input_value_reg[3][16]  ( .D(data_in[16]), .E(n354), .CP(clk), .Q(
        \input_value[3][16] ) );
  EDFQD1 \input_value_reg[3][15]  ( .D(data_in[15]), .E(n354), .CP(clk), .Q(
        \input_value[3][15] ) );
  EDFQD1 \input_value_reg[3][14]  ( .D(data_in[14]), .E(n354), .CP(clk), .Q(
        \input_value[3][14] ) );
  EDFQD1 \input_value_reg[3][13]  ( .D(data_in[13]), .E(n354), .CP(clk), .Q(
        \input_value[3][13] ) );
  EDFQD1 \input_value_reg[3][12]  ( .D(data_in[12]), .E(n353), .CP(clk), .Q(
        \input_value[3][12] ) );
  EDFQD1 \input_value_reg[3][11]  ( .D(data_in[11]), .E(n353), .CP(clk), .Q(
        \input_value[3][11] ) );
  EDFQD1 \input_value_reg[3][10]  ( .D(data_in[10]), .E(n353), .CP(clk), .Q(
        \input_value[3][10] ) );
  EDFQD1 \input_value_reg[3][9]  ( .D(data_in[9]), .E(n353), .CP(clk), .Q(
        \input_value[3][9] ) );
  EDFQD1 \input_value_reg[3][8]  ( .D(data_in[8]), .E(n353), .CP(clk), .Q(
        \input_value[3][8] ) );
  EDFQD1 \input_value_reg[3][7]  ( .D(data_in[7]), .E(n353), .CP(clk), .Q(
        \input_value[3][7] ) );
  EDFQD1 \input_value_reg[3][6]  ( .D(data_in[6]), .E(n353), .CP(clk), .Q(
        \input_value[3][6] ) );
  EDFQD1 \input_value_reg[3][5]  ( .D(data_in[5]), .E(n353), .CP(clk), .Q(
        \input_value[3][5] ) );
  EDFQD1 \input_value_reg[3][4]  ( .D(data_in[4]), .E(n353), .CP(clk), .Q(
        \input_value[3][4] ) );
  EDFQD1 \input_value_reg[3][3]  ( .D(data_in[3]), .E(n353), .CP(clk), .Q(
        \input_value[3][3] ) );
  EDFQD1 \input_value_reg[3][2]  ( .D(data_in[2]), .E(n353), .CP(clk), .Q(
        \input_value[3][2] ) );
  EDFQD1 \input_value_reg[3][1]  ( .D(data_in[1]), .E(n353), .CP(clk), .Q(
        \input_value[3][1] ) );
  EDFQD1 \input_value_reg[3][0]  ( .D(data_in[0]), .E(n353), .CP(clk), .Q(
        \input_value[3][0] ) );
  EDFQD1 \input_weight_reg[3][99]  ( .D(data_in[99]), .E(n482), .CP(clk), .Q(
        \input_weight[3][99] ) );
  EDFQD1 \input_weight_reg[3][100]  ( .D(data_in[100]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][100] ) );
  EDFQD1 \input_weight_reg[3][101]  ( .D(data_in[101]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][101] ) );
  EDFQD1 \input_weight_reg[3][102]  ( .D(data_in[102]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][102] ) );
  EDFQD1 \input_weight_reg[3][103]  ( .D(data_in[103]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][103] ) );
  EDFQD1 \input_weight_reg[3][104]  ( .D(data_in[104]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][104] ) );
  EDFQD1 \input_weight_reg[3][105]  ( .D(data_in[105]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][105] ) );
  EDFQD1 \input_weight_reg[3][106]  ( .D(data_in[106]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][106] ) );
  EDFQD1 \input_weight_reg[3][107]  ( .D(data_in[107]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][107] ) );
  EDFQD1 \input_weight_reg[3][108]  ( .D(data_in[108]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][108] ) );
  EDFQD1 \input_weight_reg[3][109]  ( .D(data_in[109]), .E(n482), .CP(clk), 
        .Q(\input_weight[3][109] ) );
  EDFQD1 \input_weight_reg[3][110]  ( .D(data_in[110]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][110] ) );
  EDFQD1 \input_weight_reg[3][111]  ( .D(data_in[111]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][111] ) );
  EDFQD1 \input_weight_reg[3][112]  ( .D(data_in[112]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][112] ) );
  EDFQD1 \input_weight_reg[3][113]  ( .D(data_in[113]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][113] ) );
  EDFQD1 \input_weight_reg[3][114]  ( .D(data_in[114]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][114] ) );
  EDFQD1 \input_weight_reg[3][115]  ( .D(data_in[115]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][115] ) );
  EDFQD1 \input_weight_reg[3][116]  ( .D(data_in[116]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][116] ) );
  EDFQD1 \input_weight_reg[3][117]  ( .D(data_in[117]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][117] ) );
  EDFQD1 \input_weight_reg[3][118]  ( .D(data_in[118]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][118] ) );
  EDFQD1 \input_weight_reg[3][119]  ( .D(data_in[119]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][119] ) );
  EDFQD1 \input_weight_reg[3][120]  ( .D(data_in[120]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][120] ) );
  EDFQD1 \input_weight_reg[3][121]  ( .D(data_in[121]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][121] ) );
  EDFQD1 \input_weight_reg[3][122]  ( .D(data_in[122]), .E(n481), .CP(clk), 
        .Q(\input_weight[3][122] ) );
  EDFQD1 \input_weight_reg[3][123]  ( .D(data_in[123]), .E(n480), .CP(clk), 
        .Q(\input_weight[3][123] ) );
  EDFQD1 \input_weight_reg[3][124]  ( .D(data_in[124]), .E(n480), .CP(clk), 
        .Q(\input_weight[3][124] ) );
  EDFQD1 \input_weight_reg[3][125]  ( .D(data_in[125]), .E(n480), .CP(clk), 
        .Q(\input_weight[3][125] ) );
  EDFQD1 \input_weight_reg[3][126]  ( .D(data_in[126]), .E(n480), .CP(clk), 
        .Q(\input_weight[3][126] ) );
  EDFQD1 \input_weight_reg[3][127]  ( .D(data_in[127]), .E(n480), .CP(clk), 
        .Q(\input_weight[3][127] ) );
  EDFQD1 \input_weight_reg[3][98]  ( .D(data_in[98]), .E(n480), .CP(clk), .Q(
        \input_weight[3][98] ) );
  EDFQD1 \input_weight_reg[3][97]  ( .D(data_in[97]), .E(n480), .CP(clk), .Q(
        \input_weight[3][97] ) );
  EDFQD1 \input_weight_reg[3][96]  ( .D(data_in[96]), .E(n480), .CP(clk), .Q(
        \input_weight[3][96] ) );
  EDFQD1 \input_weight_reg[3][95]  ( .D(data_in[95]), .E(n480), .CP(clk), .Q(
        \input_weight[3][95] ) );
  EDFQD1 \input_weight_reg[3][94]  ( .D(data_in[94]), .E(n480), .CP(clk), .Q(
        \input_weight[3][94] ) );
  EDFQD1 \input_weight_reg[3][93]  ( .D(data_in[93]), .E(n480), .CP(clk), .Q(
        \input_weight[3][93] ) );
  EDFQD1 \input_weight_reg[3][92]  ( .D(data_in[92]), .E(n480), .CP(clk), .Q(
        \input_weight[3][92] ) );
  EDFQD1 \input_weight_reg[3][91]  ( .D(data_in[91]), .E(n480), .CP(clk), .Q(
        \input_weight[3][91] ) );
  EDFQD1 \input_weight_reg[3][90]  ( .D(data_in[90]), .E(n479), .CP(clk), .Q(
        \input_weight[3][90] ) );
  EDFQD1 \input_weight_reg[3][89]  ( .D(data_in[89]), .E(n479), .CP(clk), .Q(
        \input_weight[3][89] ) );
  EDFQD1 \input_weight_reg[3][88]  ( .D(data_in[88]), .E(n479), .CP(clk), .Q(
        \input_weight[3][88] ) );
  EDFQD1 \input_weight_reg[3][87]  ( .D(data_in[87]), .E(n479), .CP(clk), .Q(
        \input_weight[3][87] ) );
  EDFQD1 \input_weight_reg[3][86]  ( .D(data_in[86]), .E(n479), .CP(clk), .Q(
        \input_weight[3][86] ) );
  EDFQD1 \input_weight_reg[3][85]  ( .D(data_in[85]), .E(n479), .CP(clk), .Q(
        \input_weight[3][85] ) );
  EDFQD1 \input_weight_reg[3][84]  ( .D(data_in[84]), .E(n479), .CP(clk), .Q(
        \input_weight[3][84] ) );
  EDFQD1 \input_weight_reg[3][83]  ( .D(data_in[83]), .E(n479), .CP(clk), .Q(
        \input_weight[3][83] ) );
  EDFQD1 \input_weight_reg[3][82]  ( .D(data_in[82]), .E(n479), .CP(clk), .Q(
        \input_weight[3][82] ) );
  EDFQD1 \input_weight_reg[3][81]  ( .D(data_in[81]), .E(n479), .CP(clk), .Q(
        \input_weight[3][81] ) );
  EDFQD1 \input_weight_reg[3][80]  ( .D(data_in[80]), .E(n479), .CP(clk), .Q(
        \input_weight[3][80] ) );
  EDFQD1 \input_weight_reg[3][79]  ( .D(data_in[79]), .E(n479), .CP(clk), .Q(
        \input_weight[3][79] ) );
  EDFQD1 \input_weight_reg[3][78]  ( .D(data_in[78]), .E(n479), .CP(clk), .Q(
        \input_weight[3][78] ) );
  EDFQD1 \input_weight_reg[3][77]  ( .D(data_in[77]), .E(n478), .CP(clk), .Q(
        \input_weight[3][77] ) );
  EDFQD1 \input_weight_reg[3][76]  ( .D(data_in[76]), .E(n478), .CP(clk), .Q(
        \input_weight[3][76] ) );
  EDFQD1 \input_weight_reg[3][75]  ( .D(data_in[75]), .E(n478), .CP(clk), .Q(
        \input_weight[3][75] ) );
  EDFQD1 \input_weight_reg[3][74]  ( .D(data_in[74]), .E(n478), .CP(clk), .Q(
        \input_weight[3][74] ) );
  EDFQD1 \input_weight_reg[3][73]  ( .D(data_in[73]), .E(n478), .CP(clk), .Q(
        \input_weight[3][73] ) );
  EDFQD1 \input_weight_reg[3][72]  ( .D(data_in[72]), .E(n478), .CP(clk), .Q(
        \input_weight[3][72] ) );
  EDFQD1 \input_weight_reg[3][71]  ( .D(data_in[71]), .E(n478), .CP(clk), .Q(
        \input_weight[3][71] ) );
  EDFQD1 \input_weight_reg[3][70]  ( .D(data_in[70]), .E(n478), .CP(clk), .Q(
        \input_weight[3][70] ) );
  EDFQD1 \input_weight_reg[3][69]  ( .D(data_in[69]), .E(n478), .CP(clk), .Q(
        \input_weight[3][69] ) );
  EDFQD1 \input_weight_reg[3][68]  ( .D(data_in[68]), .E(n478), .CP(clk), .Q(
        \input_weight[3][68] ) );
  EDFQD1 \input_weight_reg[3][67]  ( .D(data_in[67]), .E(n478), .CP(clk), .Q(
        \input_weight[3][67] ) );
  EDFQD1 \input_weight_reg[3][66]  ( .D(data_in[66]), .E(n478), .CP(clk), .Q(
        \input_weight[3][66] ) );
  EDFQD1 \input_weight_reg[3][65]  ( .D(data_in[65]), .E(n478), .CP(clk), .Q(
        \input_weight[3][65] ) );
  EDFQD1 \input_weight_reg[3][64]  ( .D(data_in[64]), .E(n477), .CP(clk), .Q(
        \input_weight[3][64] ) );
  EDFQD1 \input_weight_reg[3][63]  ( .D(data_in[63]), .E(n477), .CP(clk), .Q(
        \input_weight[3][63] ) );
  EDFQD1 \input_weight_reg[3][62]  ( .D(data_in[62]), .E(n477), .CP(clk), .Q(
        \input_weight[3][62] ) );
  EDFQD1 \input_weight_reg[3][61]  ( .D(data_in[61]), .E(n477), .CP(clk), .Q(
        \input_weight[3][61] ) );
  EDFQD1 \input_weight_reg[3][60]  ( .D(data_in[60]), .E(n477), .CP(clk), .Q(
        \input_weight[3][60] ) );
  EDFQD1 \input_weight_reg[3][59]  ( .D(data_in[59]), .E(n477), .CP(clk), .Q(
        \input_weight[3][59] ) );
  EDFQD1 \input_weight_reg[3][58]  ( .D(data_in[58]), .E(n477), .CP(clk), .Q(
        \input_weight[3][58] ) );
  EDFQD1 \input_weight_reg[3][57]  ( .D(data_in[57]), .E(n477), .CP(clk), .Q(
        \input_weight[3][57] ) );
  EDFQD1 \input_weight_reg[3][56]  ( .D(data_in[56]), .E(n477), .CP(clk), .Q(
        \input_weight[3][56] ) );
  EDFQD1 \input_weight_reg[3][55]  ( .D(data_in[55]), .E(n477), .CP(clk), .Q(
        \input_weight[3][55] ) );
  EDFQD1 \input_weight_reg[3][54]  ( .D(data_in[54]), .E(n477), .CP(clk), .Q(
        \input_weight[3][54] ) );
  EDFQD1 \input_weight_reg[3][53]  ( .D(data_in[53]), .E(n477), .CP(clk), .Q(
        \input_weight[3][53] ) );
  EDFQD1 \input_weight_reg[3][52]  ( .D(data_in[52]), .E(n477), .CP(clk), .Q(
        \input_weight[3][52] ) );
  EDFQD1 \input_weight_reg[3][51]  ( .D(data_in[51]), .E(n476), .CP(clk), .Q(
        \input_weight[3][51] ) );
  EDFQD1 \input_weight_reg[3][50]  ( .D(data_in[50]), .E(n476), .CP(clk), .Q(
        \input_weight[3][50] ) );
  EDFQD1 \input_weight_reg[3][49]  ( .D(data_in[49]), .E(n476), .CP(clk), .Q(
        \input_weight[3][49] ) );
  EDFQD1 \input_weight_reg[3][48]  ( .D(data_in[48]), .E(n476), .CP(clk), .Q(
        \input_weight[3][48] ) );
  EDFQD1 \input_weight_reg[3][47]  ( .D(data_in[47]), .E(n476), .CP(clk), .Q(
        \input_weight[3][47] ) );
  EDFQD1 \input_weight_reg[3][46]  ( .D(data_in[46]), .E(n476), .CP(clk), .Q(
        \input_weight[3][46] ) );
  EDFQD1 \input_weight_reg[3][45]  ( .D(data_in[45]), .E(n476), .CP(clk), .Q(
        \input_weight[3][45] ) );
  EDFQD1 \input_weight_reg[3][44]  ( .D(data_in[44]), .E(n476), .CP(clk), .Q(
        \input_weight[3][44] ) );
  EDFQD1 \input_weight_reg[3][43]  ( .D(data_in[43]), .E(n476), .CP(clk), .Q(
        \input_weight[3][43] ) );
  EDFQD1 \input_weight_reg[3][42]  ( .D(data_in[42]), .E(n476), .CP(clk), .Q(
        \input_weight[3][42] ) );
  EDFQD1 \input_weight_reg[3][41]  ( .D(data_in[41]), .E(n476), .CP(clk), .Q(
        \input_weight[3][41] ) );
  EDFQD1 \input_weight_reg[3][40]  ( .D(data_in[40]), .E(n476), .CP(clk), .Q(
        \input_weight[3][40] ) );
  EDFQD1 \input_weight_reg[3][39]  ( .D(data_in[39]), .E(n476), .CP(clk), .Q(
        \input_weight[3][39] ) );
  EDFQD1 \input_weight_reg[3][38]  ( .D(data_in[38]), .E(n475), .CP(clk), .Q(
        \input_weight[3][38] ) );
  EDFQD1 \input_weight_reg[3][37]  ( .D(data_in[37]), .E(n475), .CP(clk), .Q(
        \input_weight[3][37] ) );
  EDFQD1 \input_weight_reg[3][36]  ( .D(data_in[36]), .E(n475), .CP(clk), .Q(
        \input_weight[3][36] ) );
  EDFQD1 \input_weight_reg[3][35]  ( .D(data_in[35]), .E(n475), .CP(clk), .Q(
        \input_weight[3][35] ) );
  EDFQD1 \input_weight_reg[3][34]  ( .D(data_in[34]), .E(n475), .CP(clk), .Q(
        \input_weight[3][34] ) );
  EDFQD1 \input_weight_reg[3][33]  ( .D(data_in[33]), .E(n475), .CP(clk), .Q(
        \input_weight[3][33] ) );
  EDFQD1 \input_weight_reg[3][32]  ( .D(data_in[32]), .E(n475), .CP(clk), .Q(
        \input_weight[3][32] ) );
  EDFQD1 \input_weight_reg[3][31]  ( .D(data_in[31]), .E(n475), .CP(clk), .Q(
        \input_weight[3][31] ) );
  EDFQD1 \input_weight_reg[3][30]  ( .D(data_in[30]), .E(n475), .CP(clk), .Q(
        \input_weight[3][30] ) );
  EDFQD1 \input_weight_reg[3][29]  ( .D(data_in[29]), .E(n475), .CP(clk), .Q(
        \input_weight[3][29] ) );
  EDFQD1 \input_weight_reg[3][28]  ( .D(data_in[28]), .E(n475), .CP(clk), .Q(
        \input_weight[3][28] ) );
  EDFQD1 \input_weight_reg[3][27]  ( .D(data_in[27]), .E(n475), .CP(clk), .Q(
        \input_weight[3][27] ) );
  EDFQD1 \input_weight_reg[3][26]  ( .D(data_in[26]), .E(n475), .CP(clk), .Q(
        \input_weight[3][26] ) );
  EDFQD1 \input_weight_reg[3][25]  ( .D(data_in[25]), .E(n474), .CP(clk), .Q(
        \input_weight[3][25] ) );
  EDFQD1 \input_weight_reg[3][24]  ( .D(data_in[24]), .E(n474), .CP(clk), .Q(
        \input_weight[3][24] ) );
  EDFQD1 \input_weight_reg[3][23]  ( .D(data_in[23]), .E(n474), .CP(clk), .Q(
        \input_weight[3][23] ) );
  EDFQD1 \input_weight_reg[3][22]  ( .D(data_in[22]), .E(n474), .CP(clk), .Q(
        \input_weight[3][22] ) );
  EDFQD1 \input_weight_reg[3][21]  ( .D(data_in[21]), .E(n474), .CP(clk), .Q(
        \input_weight[3][21] ) );
  EDFQD1 \input_weight_reg[3][20]  ( .D(data_in[20]), .E(n474), .CP(clk), .Q(
        \input_weight[3][20] ) );
  EDFQD1 \input_weight_reg[3][19]  ( .D(data_in[19]), .E(n474), .CP(clk), .Q(
        \input_weight[3][19] ) );
  EDFQD1 \input_weight_reg[3][18]  ( .D(data_in[18]), .E(n474), .CP(clk), .Q(
        \input_weight[3][18] ) );
  EDFQD1 \input_weight_reg[3][17]  ( .D(data_in[17]), .E(n474), .CP(clk), .Q(
        \input_weight[3][17] ) );
  EDFQD1 \input_weight_reg[3][16]  ( .D(data_in[16]), .E(n474), .CP(clk), .Q(
        \input_weight[3][16] ) );
  EDFQD1 \input_weight_reg[3][15]  ( .D(data_in[15]), .E(n474), .CP(clk), .Q(
        \input_weight[3][15] ) );
  EDFQD1 \input_weight_reg[3][14]  ( .D(data_in[14]), .E(n474), .CP(clk), .Q(
        \input_weight[3][14] ) );
  EDFQD1 \input_weight_reg[3][13]  ( .D(data_in[13]), .E(n474), .CP(clk), .Q(
        \input_weight[3][13] ) );
  EDFQD1 \input_weight_reg[3][12]  ( .D(data_in[12]), .E(n473), .CP(clk), .Q(
        \input_weight[3][12] ) );
  EDFQD1 \input_weight_reg[3][11]  ( .D(data_in[11]), .E(n473), .CP(clk), .Q(
        \input_weight[3][11] ) );
  EDFQD1 \input_weight_reg[3][10]  ( .D(data_in[10]), .E(n473), .CP(clk), .Q(
        \input_weight[3][10] ) );
  EDFQD1 \input_weight_reg[3][9]  ( .D(data_in[9]), .E(n473), .CP(clk), .Q(
        \input_weight[3][9] ) );
  EDFQD1 \input_weight_reg[3][8]  ( .D(data_in[8]), .E(n473), .CP(clk), .Q(
        \input_weight[3][8] ) );
  EDFQD1 \input_weight_reg[3][7]  ( .D(data_in[7]), .E(n473), .CP(clk), .Q(
        \input_weight[3][7] ) );
  EDFQD1 \input_weight_reg[3][6]  ( .D(data_in[6]), .E(n473), .CP(clk), .Q(
        \input_weight[3][6] ) );
  EDFQD1 \input_weight_reg[3][5]  ( .D(data_in[5]), .E(n473), .CP(clk), .Q(
        \input_weight[3][5] ) );
  EDFQD1 \input_weight_reg[3][4]  ( .D(data_in[4]), .E(n473), .CP(clk), .Q(
        \input_weight[3][4] ) );
  EDFQD1 \input_weight_reg[3][3]  ( .D(data_in[3]), .E(n473), .CP(clk), .Q(
        \input_weight[3][3] ) );
  EDFQD1 \input_weight_reg[3][2]  ( .D(data_in[2]), .E(n473), .CP(clk), .Q(
        \input_weight[3][2] ) );
  EDFQD1 \input_weight_reg[3][1]  ( .D(data_in[1]), .E(n473), .CP(clk), .Q(
        \input_weight[3][1] ) );
  EDFQD1 \input_weight_reg[3][0]  ( .D(data_in[0]), .E(n473), .CP(clk), .Q(
        \input_weight[3][0] ) );
  EDFQD1 \input_value_reg[4][99]  ( .D(data_in[99]), .E(n347), .CP(clk), .Q(
        \input_value[4][99] ) );
  EDFQD1 \input_value_reg[4][100]  ( .D(data_in[100]), .E(n347), .CP(clk), .Q(
        \input_value[4][100] ) );
  EDFQD1 \input_value_reg[4][101]  ( .D(data_in[101]), .E(n347), .CP(clk), .Q(
        \input_value[4][101] ) );
  EDFQD1 \input_value_reg[4][102]  ( .D(data_in[102]), .E(n347), .CP(clk), .Q(
        \input_value[4][102] ) );
  EDFQD1 \input_value_reg[4][103]  ( .D(data_in[103]), .E(n347), .CP(clk), .Q(
        \input_value[4][103] ) );
  EDFQD1 \input_value_reg[4][104]  ( .D(data_in[104]), .E(n347), .CP(clk), .Q(
        \input_value[4][104] ) );
  EDFQD1 \input_value_reg[4][105]  ( .D(data_in[105]), .E(n347), .CP(clk), .Q(
        \input_value[4][105] ) );
  EDFQD1 \input_value_reg[4][106]  ( .D(data_in[106]), .E(n347), .CP(clk), .Q(
        \input_value[4][106] ) );
  EDFQD1 \input_value_reg[4][107]  ( .D(data_in[107]), .E(n347), .CP(clk), .Q(
        \input_value[4][107] ) );
  EDFQD1 \input_value_reg[4][108]  ( .D(data_in[108]), .E(n347), .CP(clk), .Q(
        \input_value[4][108] ) );
  EDFQD1 \input_value_reg[4][109]  ( .D(data_in[109]), .E(n347), .CP(clk), .Q(
        \input_value[4][109] ) );
  EDFQD1 \input_value_reg[4][110]  ( .D(data_in[110]), .E(n346), .CP(clk), .Q(
        \input_value[4][110] ) );
  EDFQD1 \input_value_reg[4][111]  ( .D(data_in[111]), .E(n346), .CP(clk), .Q(
        \input_value[4][111] ) );
  EDFQD1 \input_value_reg[4][112]  ( .D(data_in[112]), .E(n346), .CP(clk), .Q(
        \input_value[4][112] ) );
  EDFQD1 \input_value_reg[4][113]  ( .D(data_in[113]), .E(n346), .CP(clk), .Q(
        \input_value[4][113] ) );
  EDFQD1 \input_value_reg[4][114]  ( .D(data_in[114]), .E(n346), .CP(clk), .Q(
        \input_value[4][114] ) );
  EDFQD1 \input_value_reg[4][115]  ( .D(data_in[115]), .E(n346), .CP(clk), .Q(
        \input_value[4][115] ) );
  EDFQD1 \input_value_reg[4][116]  ( .D(data_in[116]), .E(n346), .CP(clk), .Q(
        \input_value[4][116] ) );
  EDFQD1 \input_value_reg[4][117]  ( .D(data_in[117]), .E(n346), .CP(clk), .Q(
        \input_value[4][117] ) );
  EDFQD1 \input_value_reg[4][118]  ( .D(data_in[118]), .E(n346), .CP(clk), .Q(
        \input_value[4][118] ) );
  EDFQD1 \input_value_reg[4][119]  ( .D(data_in[119]), .E(n346), .CP(clk), .Q(
        \input_value[4][119] ) );
  EDFQD1 \input_value_reg[4][120]  ( .D(data_in[120]), .E(n346), .CP(clk), .Q(
        \input_value[4][120] ) );
  EDFQD1 \input_value_reg[4][121]  ( .D(data_in[121]), .E(n346), .CP(clk), .Q(
        \input_value[4][121] ) );
  EDFQD1 \input_value_reg[4][122]  ( .D(data_in[122]), .E(n346), .CP(clk), .Q(
        \input_value[4][122] ) );
  EDFQD1 \input_value_reg[4][123]  ( .D(data_in[123]), .E(n345), .CP(clk), .Q(
        \input_value[4][123] ) );
  EDFQD1 \input_value_reg[4][124]  ( .D(data_in[124]), .E(n345), .CP(clk), .Q(
        \input_value[4][124] ) );
  EDFQD1 \input_value_reg[4][125]  ( .D(data_in[125]), .E(n345), .CP(clk), .Q(
        \input_value[4][125] ) );
  EDFQD1 \input_value_reg[4][126]  ( .D(data_in[126]), .E(n345), .CP(clk), .Q(
        \input_value[4][126] ) );
  EDFQD1 \input_value_reg[4][127]  ( .D(data_in[127]), .E(n345), .CP(clk), .Q(
        \input_value[4][127] ) );
  EDFQD1 \input_value_reg[4][98]  ( .D(data_in[98]), .E(n345), .CP(clk), .Q(
        \input_value[4][98] ) );
  EDFQD1 \input_value_reg[4][97]  ( .D(data_in[97]), .E(n345), .CP(clk), .Q(
        \input_value[4][97] ) );
  EDFQD1 \input_value_reg[4][96]  ( .D(data_in[96]), .E(n345), .CP(clk), .Q(
        \input_value[4][96] ) );
  EDFQD1 \input_value_reg[4][95]  ( .D(data_in[95]), .E(n345), .CP(clk), .Q(
        \input_value[4][95] ) );
  EDFQD1 \input_value_reg[4][94]  ( .D(data_in[94]), .E(n345), .CP(clk), .Q(
        \input_value[4][94] ) );
  EDFQD1 \input_value_reg[4][93]  ( .D(data_in[93]), .E(n345), .CP(clk), .Q(
        \input_value[4][93] ) );
  EDFQD1 \input_value_reg[4][92]  ( .D(data_in[92]), .E(n345), .CP(clk), .Q(
        \input_value[4][92] ) );
  EDFQD1 \input_value_reg[4][91]  ( .D(data_in[91]), .E(n345), .CP(clk), .Q(
        \input_value[4][91] ) );
  EDFQD1 \input_value_reg[4][90]  ( .D(data_in[90]), .E(n344), .CP(clk), .Q(
        \input_value[4][90] ) );
  EDFQD1 \input_value_reg[4][89]  ( .D(data_in[89]), .E(n344), .CP(clk), .Q(
        \input_value[4][89] ) );
  EDFQD1 \input_value_reg[4][88]  ( .D(data_in[88]), .E(n344), .CP(clk), .Q(
        \input_value[4][88] ) );
  EDFQD1 \input_value_reg[4][87]  ( .D(data_in[87]), .E(n344), .CP(clk), .Q(
        \input_value[4][87] ) );
  EDFQD1 \input_value_reg[4][86]  ( .D(data_in[86]), .E(n344), .CP(clk), .Q(
        \input_value[4][86] ) );
  EDFQD1 \input_value_reg[4][85]  ( .D(data_in[85]), .E(n344), .CP(clk), .Q(
        \input_value[4][85] ) );
  EDFQD1 \input_value_reg[4][84]  ( .D(data_in[84]), .E(n344), .CP(clk), .Q(
        \input_value[4][84] ) );
  EDFQD1 \input_value_reg[4][83]  ( .D(data_in[83]), .E(n344), .CP(clk), .Q(
        \input_value[4][83] ) );
  EDFQD1 \input_value_reg[4][82]  ( .D(data_in[82]), .E(n344), .CP(clk), .Q(
        \input_value[4][82] ) );
  EDFQD1 \input_value_reg[4][81]  ( .D(data_in[81]), .E(n344), .CP(clk), .Q(
        \input_value[4][81] ) );
  EDFQD1 \input_value_reg[4][80]  ( .D(data_in[80]), .E(n344), .CP(clk), .Q(
        \input_value[4][80] ) );
  EDFQD1 \input_value_reg[4][79]  ( .D(data_in[79]), .E(n344), .CP(clk), .Q(
        \input_value[4][79] ) );
  EDFQD1 \input_value_reg[4][78]  ( .D(data_in[78]), .E(n344), .CP(clk), .Q(
        \input_value[4][78] ) );
  EDFQD1 \input_value_reg[4][77]  ( .D(data_in[77]), .E(n343), .CP(clk), .Q(
        \input_value[4][77] ) );
  EDFQD1 \input_value_reg[4][76]  ( .D(data_in[76]), .E(n343), .CP(clk), .Q(
        \input_value[4][76] ) );
  EDFQD1 \input_value_reg[4][75]  ( .D(data_in[75]), .E(n343), .CP(clk), .Q(
        \input_value[4][75] ) );
  EDFQD1 \input_value_reg[4][74]  ( .D(data_in[74]), .E(n343), .CP(clk), .Q(
        \input_value[4][74] ) );
  EDFQD1 \input_value_reg[4][73]  ( .D(data_in[73]), .E(n343), .CP(clk), .Q(
        \input_value[4][73] ) );
  EDFQD1 \input_value_reg[4][72]  ( .D(data_in[72]), .E(n343), .CP(clk), .Q(
        \input_value[4][72] ) );
  EDFQD1 \input_value_reg[4][71]  ( .D(data_in[71]), .E(n343), .CP(clk), .Q(
        \input_value[4][71] ) );
  EDFQD1 \input_value_reg[4][70]  ( .D(data_in[70]), .E(n343), .CP(clk), .Q(
        \input_value[4][70] ) );
  EDFQD1 \input_value_reg[4][69]  ( .D(data_in[69]), .E(n343), .CP(clk), .Q(
        \input_value[4][69] ) );
  EDFQD1 \input_value_reg[4][68]  ( .D(data_in[68]), .E(n343), .CP(clk), .Q(
        \input_value[4][68] ) );
  EDFQD1 \input_value_reg[4][67]  ( .D(data_in[67]), .E(n343), .CP(clk), .Q(
        \input_value[4][67] ) );
  EDFQD1 \input_value_reg[4][66]  ( .D(data_in[66]), .E(n343), .CP(clk), .Q(
        \input_value[4][66] ) );
  EDFQD1 \input_value_reg[4][65]  ( .D(data_in[65]), .E(n343), .CP(clk), .Q(
        \input_value[4][65] ) );
  EDFQD1 \input_value_reg[4][64]  ( .D(data_in[64]), .E(n342), .CP(clk), .Q(
        \input_value[4][64] ) );
  EDFQD1 \input_value_reg[4][63]  ( .D(data_in[63]), .E(n342), .CP(clk), .Q(
        \input_value[4][63] ) );
  EDFQD1 \input_value_reg[4][62]  ( .D(data_in[62]), .E(n342), .CP(clk), .Q(
        \input_value[4][62] ) );
  EDFQD1 \input_value_reg[4][61]  ( .D(data_in[61]), .E(n342), .CP(clk), .Q(
        \input_value[4][61] ) );
  EDFQD1 \input_value_reg[4][60]  ( .D(data_in[60]), .E(n342), .CP(clk), .Q(
        \input_value[4][60] ) );
  EDFQD1 \input_value_reg[4][59]  ( .D(data_in[59]), .E(n342), .CP(clk), .Q(
        \input_value[4][59] ) );
  EDFQD1 \input_value_reg[4][58]  ( .D(data_in[58]), .E(n342), .CP(clk), .Q(
        \input_value[4][58] ) );
  EDFQD1 \input_value_reg[4][57]  ( .D(data_in[57]), .E(n342), .CP(clk), .Q(
        \input_value[4][57] ) );
  EDFQD1 \input_value_reg[4][56]  ( .D(data_in[56]), .E(n342), .CP(clk), .Q(
        \input_value[4][56] ) );
  EDFQD1 \input_value_reg[4][55]  ( .D(data_in[55]), .E(n342), .CP(clk), .Q(
        \input_value[4][55] ) );
  EDFQD1 \input_value_reg[4][54]  ( .D(data_in[54]), .E(n342), .CP(clk), .Q(
        \input_value[4][54] ) );
  EDFQD1 \input_value_reg[4][53]  ( .D(data_in[53]), .E(n342), .CP(clk), .Q(
        \input_value[4][53] ) );
  EDFQD1 \input_value_reg[4][52]  ( .D(data_in[52]), .E(n342), .CP(clk), .Q(
        \input_value[4][52] ) );
  EDFQD1 \input_value_reg[4][51]  ( .D(data_in[51]), .E(n341), .CP(clk), .Q(
        \input_value[4][51] ) );
  EDFQD1 \input_value_reg[4][50]  ( .D(data_in[50]), .E(n341), .CP(clk), .Q(
        \input_value[4][50] ) );
  EDFQD1 \input_value_reg[4][49]  ( .D(data_in[49]), .E(n341), .CP(clk), .Q(
        \input_value[4][49] ) );
  EDFQD1 \input_value_reg[4][48]  ( .D(data_in[48]), .E(n341), .CP(clk), .Q(
        \input_value[4][48] ) );
  EDFQD1 \input_value_reg[4][47]  ( .D(data_in[47]), .E(n341), .CP(clk), .Q(
        \input_value[4][47] ) );
  EDFQD1 \input_value_reg[4][46]  ( .D(data_in[46]), .E(n341), .CP(clk), .Q(
        \input_value[4][46] ) );
  EDFQD1 \input_value_reg[4][45]  ( .D(data_in[45]), .E(n341), .CP(clk), .Q(
        \input_value[4][45] ) );
  EDFQD1 \input_value_reg[4][44]  ( .D(data_in[44]), .E(n341), .CP(clk), .Q(
        \input_value[4][44] ) );
  EDFQD1 \input_value_reg[4][43]  ( .D(data_in[43]), .E(n341), .CP(clk), .Q(
        \input_value[4][43] ) );
  EDFQD1 \input_value_reg[4][42]  ( .D(data_in[42]), .E(n341), .CP(clk), .Q(
        \input_value[4][42] ) );
  EDFQD1 \input_value_reg[4][41]  ( .D(data_in[41]), .E(n341), .CP(clk), .Q(
        \input_value[4][41] ) );
  EDFQD1 \input_value_reg[4][40]  ( .D(data_in[40]), .E(n341), .CP(clk), .Q(
        \input_value[4][40] ) );
  EDFQD1 \input_value_reg[4][39]  ( .D(data_in[39]), .E(n341), .CP(clk), .Q(
        \input_value[4][39] ) );
  EDFQD1 \input_value_reg[4][38]  ( .D(data_in[38]), .E(n340), .CP(clk), .Q(
        \input_value[4][38] ) );
  EDFQD1 \input_value_reg[4][37]  ( .D(data_in[37]), .E(n340), .CP(clk), .Q(
        \input_value[4][37] ) );
  EDFQD1 \input_value_reg[4][36]  ( .D(data_in[36]), .E(n340), .CP(clk), .Q(
        \input_value[4][36] ) );
  EDFQD1 \input_value_reg[4][35]  ( .D(data_in[35]), .E(n340), .CP(clk), .Q(
        \input_value[4][35] ) );
  EDFQD1 \input_value_reg[4][34]  ( .D(data_in[34]), .E(n340), .CP(clk), .Q(
        \input_value[4][34] ) );
  EDFQD1 \input_value_reg[4][33]  ( .D(data_in[33]), .E(n340), .CP(clk), .Q(
        \input_value[4][33] ) );
  EDFQD1 \input_value_reg[4][32]  ( .D(data_in[32]), .E(n340), .CP(clk), .Q(
        \input_value[4][32] ) );
  EDFQD1 \input_value_reg[4][31]  ( .D(data_in[31]), .E(n340), .CP(clk), .Q(
        \input_value[4][31] ) );
  EDFQD1 \input_value_reg[4][30]  ( .D(data_in[30]), .E(n340), .CP(clk), .Q(
        \input_value[4][30] ) );
  EDFQD1 \input_value_reg[4][29]  ( .D(data_in[29]), .E(n340), .CP(clk), .Q(
        \input_value[4][29] ) );
  EDFQD1 \input_value_reg[4][28]  ( .D(data_in[28]), .E(n340), .CP(clk), .Q(
        \input_value[4][28] ) );
  EDFQD1 \input_value_reg[4][27]  ( .D(data_in[27]), .E(n340), .CP(clk), .Q(
        \input_value[4][27] ) );
  EDFQD1 \input_value_reg[4][26]  ( .D(data_in[26]), .E(n340), .CP(clk), .Q(
        \input_value[4][26] ) );
  EDFQD1 \input_value_reg[4][25]  ( .D(data_in[25]), .E(n339), .CP(clk), .Q(
        \input_value[4][25] ) );
  EDFQD1 \input_value_reg[4][24]  ( .D(data_in[24]), .E(n339), .CP(clk), .Q(
        \input_value[4][24] ) );
  EDFQD1 \input_value_reg[4][23]  ( .D(data_in[23]), .E(n339), .CP(clk), .Q(
        \input_value[4][23] ) );
  EDFQD1 \input_value_reg[4][22]  ( .D(data_in[22]), .E(n339), .CP(clk), .Q(
        \input_value[4][22] ) );
  EDFQD1 \input_value_reg[4][21]  ( .D(data_in[21]), .E(n339), .CP(clk), .Q(
        \input_value[4][21] ) );
  EDFQD1 \input_value_reg[4][20]  ( .D(data_in[20]), .E(n339), .CP(clk), .Q(
        \input_value[4][20] ) );
  EDFQD1 \input_value_reg[4][19]  ( .D(data_in[19]), .E(n339), .CP(clk), .Q(
        \input_value[4][19] ) );
  EDFQD1 \input_value_reg[4][18]  ( .D(data_in[18]), .E(n339), .CP(clk), .Q(
        \input_value[4][18] ) );
  EDFQD1 \input_value_reg[4][17]  ( .D(data_in[17]), .E(n339), .CP(clk), .Q(
        \input_value[4][17] ) );
  EDFQD1 \input_value_reg[4][16]  ( .D(data_in[16]), .E(n339), .CP(clk), .Q(
        \input_value[4][16] ) );
  EDFQD1 \input_value_reg[4][15]  ( .D(data_in[15]), .E(n339), .CP(clk), .Q(
        \input_value[4][15] ) );
  EDFQD1 \input_value_reg[4][14]  ( .D(data_in[14]), .E(n339), .CP(clk), .Q(
        \input_value[4][14] ) );
  EDFQD1 \input_value_reg[4][13]  ( .D(data_in[13]), .E(n339), .CP(clk), .Q(
        \input_value[4][13] ) );
  EDFQD1 \input_value_reg[4][12]  ( .D(data_in[12]), .E(n338), .CP(clk), .Q(
        \input_value[4][12] ) );
  EDFQD1 \input_value_reg[4][11]  ( .D(data_in[11]), .E(n338), .CP(clk), .Q(
        \input_value[4][11] ) );
  EDFQD1 \input_value_reg[4][10]  ( .D(data_in[10]), .E(n338), .CP(clk), .Q(
        \input_value[4][10] ) );
  EDFQD1 \input_value_reg[4][9]  ( .D(data_in[9]), .E(n338), .CP(clk), .Q(
        \input_value[4][9] ) );
  EDFQD1 \input_value_reg[4][8]  ( .D(data_in[8]), .E(n338), .CP(clk), .Q(
        \input_value[4][8] ) );
  EDFQD1 \input_value_reg[4][7]  ( .D(data_in[7]), .E(n338), .CP(clk), .Q(
        \input_value[4][7] ) );
  EDFQD1 \input_value_reg[4][6]  ( .D(data_in[6]), .E(n338), .CP(clk), .Q(
        \input_value[4][6] ) );
  EDFQD1 \input_value_reg[4][5]  ( .D(data_in[5]), .E(n338), .CP(clk), .Q(
        \input_value[4][5] ) );
  EDFQD1 \input_value_reg[4][4]  ( .D(data_in[4]), .E(n338), .CP(clk), .Q(
        \input_value[4][4] ) );
  EDFQD1 \input_value_reg[4][3]  ( .D(data_in[3]), .E(n338), .CP(clk), .Q(
        \input_value[4][3] ) );
  EDFQD1 \input_value_reg[4][2]  ( .D(data_in[2]), .E(n338), .CP(clk), .Q(
        \input_value[4][2] ) );
  EDFQD1 \input_value_reg[4][1]  ( .D(data_in[1]), .E(n338), .CP(clk), .Q(
        \input_value[4][1] ) );
  EDFQD1 \input_value_reg[4][0]  ( .D(data_in[0]), .E(n338), .CP(clk), .Q(
        \input_value[4][0] ) );
  EDFQD1 \input_weight_reg[4][99]  ( .D(data_in[99]), .E(n467), .CP(clk), .Q(
        \input_weight[4][99] ) );
  EDFQD1 \input_weight_reg[4][100]  ( .D(data_in[100]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][100] ) );
  EDFQD1 \input_weight_reg[4][101]  ( .D(data_in[101]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][101] ) );
  EDFQD1 \input_weight_reg[4][102]  ( .D(data_in[102]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][102] ) );
  EDFQD1 \input_weight_reg[4][103]  ( .D(data_in[103]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][103] ) );
  EDFQD1 \input_weight_reg[4][104]  ( .D(data_in[104]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][104] ) );
  EDFQD1 \input_weight_reg[4][105]  ( .D(data_in[105]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][105] ) );
  EDFQD1 \input_weight_reg[4][106]  ( .D(data_in[106]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][106] ) );
  EDFQD1 \input_weight_reg[4][107]  ( .D(data_in[107]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][107] ) );
  EDFQD1 \input_weight_reg[4][108]  ( .D(data_in[108]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][108] ) );
  EDFQD1 \input_weight_reg[4][109]  ( .D(data_in[109]), .E(n467), .CP(clk), 
        .Q(\input_weight[4][109] ) );
  EDFQD1 \input_weight_reg[4][110]  ( .D(data_in[110]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][110] ) );
  EDFQD1 \input_weight_reg[4][111]  ( .D(data_in[111]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][111] ) );
  EDFQD1 \input_weight_reg[4][112]  ( .D(data_in[112]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][112] ) );
  EDFQD1 \input_weight_reg[4][113]  ( .D(data_in[113]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][113] ) );
  EDFQD1 \input_weight_reg[4][114]  ( .D(data_in[114]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][114] ) );
  EDFQD1 \input_weight_reg[4][115]  ( .D(data_in[115]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][115] ) );
  EDFQD1 \input_weight_reg[4][116]  ( .D(data_in[116]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][116] ) );
  EDFQD1 \input_weight_reg[4][117]  ( .D(data_in[117]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][117] ) );
  EDFQD1 \input_weight_reg[4][118]  ( .D(data_in[118]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][118] ) );
  EDFQD1 \input_weight_reg[4][119]  ( .D(data_in[119]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][119] ) );
  EDFQD1 \input_weight_reg[4][120]  ( .D(data_in[120]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][120] ) );
  EDFQD1 \input_weight_reg[4][121]  ( .D(data_in[121]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][121] ) );
  EDFQD1 \input_weight_reg[4][122]  ( .D(data_in[122]), .E(n466), .CP(clk), 
        .Q(\input_weight[4][122] ) );
  EDFQD1 \input_weight_reg[4][123]  ( .D(data_in[123]), .E(n465), .CP(clk), 
        .Q(\input_weight[4][123] ) );
  EDFQD1 \input_weight_reg[4][124]  ( .D(data_in[124]), .E(n465), .CP(clk), 
        .Q(\input_weight[4][124] ) );
  EDFQD1 \input_weight_reg[4][125]  ( .D(data_in[125]), .E(n465), .CP(clk), 
        .Q(\input_weight[4][125] ) );
  EDFQD1 \input_weight_reg[4][126]  ( .D(data_in[126]), .E(n465), .CP(clk), 
        .Q(\input_weight[4][126] ) );
  EDFQD1 \input_weight_reg[4][127]  ( .D(data_in[127]), .E(n465), .CP(clk), 
        .Q(\input_weight[4][127] ) );
  EDFQD1 \input_weight_reg[4][98]  ( .D(data_in[98]), .E(n465), .CP(clk), .Q(
        \input_weight[4][98] ) );
  EDFQD1 \input_weight_reg[4][97]  ( .D(data_in[97]), .E(n465), .CP(clk), .Q(
        \input_weight[4][97] ) );
  EDFQD1 \input_weight_reg[4][96]  ( .D(data_in[96]), .E(n465), .CP(clk), .Q(
        \input_weight[4][96] ) );
  EDFQD1 \input_weight_reg[4][95]  ( .D(data_in[95]), .E(n465), .CP(clk), .Q(
        \input_weight[4][95] ) );
  EDFQD1 \input_weight_reg[4][94]  ( .D(data_in[94]), .E(n465), .CP(clk), .Q(
        \input_weight[4][94] ) );
  EDFQD1 \input_weight_reg[4][93]  ( .D(data_in[93]), .E(n465), .CP(clk), .Q(
        \input_weight[4][93] ) );
  EDFQD1 \input_weight_reg[4][92]  ( .D(data_in[92]), .E(n465), .CP(clk), .Q(
        \input_weight[4][92] ) );
  EDFQD1 \input_weight_reg[4][91]  ( .D(data_in[91]), .E(n465), .CP(clk), .Q(
        \input_weight[4][91] ) );
  EDFQD1 \input_weight_reg[4][90]  ( .D(data_in[90]), .E(n464), .CP(clk), .Q(
        \input_weight[4][90] ) );
  EDFQD1 \input_weight_reg[4][89]  ( .D(data_in[89]), .E(n464), .CP(clk), .Q(
        \input_weight[4][89] ) );
  EDFQD1 \input_weight_reg[4][88]  ( .D(data_in[88]), .E(n464), .CP(clk), .Q(
        \input_weight[4][88] ) );
  EDFQD1 \input_weight_reg[4][87]  ( .D(data_in[87]), .E(n464), .CP(clk), .Q(
        \input_weight[4][87] ) );
  EDFQD1 \input_weight_reg[4][86]  ( .D(data_in[86]), .E(n464), .CP(clk), .Q(
        \input_weight[4][86] ) );
  EDFQD1 \input_weight_reg[4][85]  ( .D(data_in[85]), .E(n464), .CP(clk), .Q(
        \input_weight[4][85] ) );
  EDFQD1 \input_weight_reg[4][84]  ( .D(data_in[84]), .E(n464), .CP(clk), .Q(
        \input_weight[4][84] ) );
  EDFQD1 \input_weight_reg[4][83]  ( .D(data_in[83]), .E(n464), .CP(clk), .Q(
        \input_weight[4][83] ) );
  EDFQD1 \input_weight_reg[4][82]  ( .D(data_in[82]), .E(n464), .CP(clk), .Q(
        \input_weight[4][82] ) );
  EDFQD1 \input_weight_reg[4][81]  ( .D(data_in[81]), .E(n464), .CP(clk), .Q(
        \input_weight[4][81] ) );
  EDFQD1 \input_weight_reg[4][80]  ( .D(data_in[80]), .E(n464), .CP(clk), .Q(
        \input_weight[4][80] ) );
  EDFQD1 \input_weight_reg[4][79]  ( .D(data_in[79]), .E(n464), .CP(clk), .Q(
        \input_weight[4][79] ) );
  EDFQD1 \input_weight_reg[4][78]  ( .D(data_in[78]), .E(n464), .CP(clk), .Q(
        \input_weight[4][78] ) );
  EDFQD1 \input_weight_reg[4][77]  ( .D(data_in[77]), .E(n463), .CP(clk), .Q(
        \input_weight[4][77] ) );
  EDFQD1 \input_weight_reg[4][76]  ( .D(data_in[76]), .E(n463), .CP(clk), .Q(
        \input_weight[4][76] ) );
  EDFQD1 \input_weight_reg[4][75]  ( .D(data_in[75]), .E(n463), .CP(clk), .Q(
        \input_weight[4][75] ) );
  EDFQD1 \input_weight_reg[4][74]  ( .D(data_in[74]), .E(n463), .CP(clk), .Q(
        \input_weight[4][74] ) );
  EDFQD1 \input_weight_reg[4][73]  ( .D(data_in[73]), .E(n463), .CP(clk), .Q(
        \input_weight[4][73] ) );
  EDFQD1 \input_weight_reg[4][72]  ( .D(data_in[72]), .E(n463), .CP(clk), .Q(
        \input_weight[4][72] ) );
  EDFQD1 \input_weight_reg[4][71]  ( .D(data_in[71]), .E(n463), .CP(clk), .Q(
        \input_weight[4][71] ) );
  EDFQD1 \input_weight_reg[4][70]  ( .D(data_in[70]), .E(n463), .CP(clk), .Q(
        \input_weight[4][70] ) );
  EDFQD1 \input_weight_reg[4][69]  ( .D(data_in[69]), .E(n463), .CP(clk), .Q(
        \input_weight[4][69] ) );
  EDFQD1 \input_weight_reg[4][68]  ( .D(data_in[68]), .E(n463), .CP(clk), .Q(
        \input_weight[4][68] ) );
  EDFQD1 \input_weight_reg[4][67]  ( .D(data_in[67]), .E(n463), .CP(clk), .Q(
        \input_weight[4][67] ) );
  EDFQD1 \input_weight_reg[4][66]  ( .D(data_in[66]), .E(n463), .CP(clk), .Q(
        \input_weight[4][66] ) );
  EDFQD1 \input_weight_reg[4][65]  ( .D(data_in[65]), .E(n463), .CP(clk), .Q(
        \input_weight[4][65] ) );
  EDFQD1 \input_weight_reg[4][64]  ( .D(data_in[64]), .E(n462), .CP(clk), .Q(
        \input_weight[4][64] ) );
  EDFQD1 \input_weight_reg[4][63]  ( .D(data_in[63]), .E(n462), .CP(clk), .Q(
        \input_weight[4][63] ) );
  EDFQD1 \input_weight_reg[4][62]  ( .D(data_in[62]), .E(n462), .CP(clk), .Q(
        \input_weight[4][62] ) );
  EDFQD1 \input_weight_reg[4][61]  ( .D(data_in[61]), .E(n462), .CP(clk), .Q(
        \input_weight[4][61] ) );
  EDFQD1 \input_weight_reg[4][60]  ( .D(data_in[60]), .E(n462), .CP(clk), .Q(
        \input_weight[4][60] ) );
  EDFQD1 \input_weight_reg[4][59]  ( .D(data_in[59]), .E(n462), .CP(clk), .Q(
        \input_weight[4][59] ) );
  EDFQD1 \input_weight_reg[4][58]  ( .D(data_in[58]), .E(n462), .CP(clk), .Q(
        \input_weight[4][58] ) );
  EDFQD1 \input_weight_reg[4][57]  ( .D(data_in[57]), .E(n462), .CP(clk), .Q(
        \input_weight[4][57] ) );
  EDFQD1 \input_weight_reg[4][56]  ( .D(data_in[56]), .E(n462), .CP(clk), .Q(
        \input_weight[4][56] ) );
  EDFQD1 \input_weight_reg[4][55]  ( .D(data_in[55]), .E(n462), .CP(clk), .Q(
        \input_weight[4][55] ) );
  EDFQD1 \input_weight_reg[4][54]  ( .D(data_in[54]), .E(n462), .CP(clk), .Q(
        \input_weight[4][54] ) );
  EDFQD1 \input_weight_reg[4][53]  ( .D(data_in[53]), .E(n462), .CP(clk), .Q(
        \input_weight[4][53] ) );
  EDFQD1 \input_weight_reg[4][52]  ( .D(data_in[52]), .E(n462), .CP(clk), .Q(
        \input_weight[4][52] ) );
  EDFQD1 \input_weight_reg[4][51]  ( .D(data_in[51]), .E(n461), .CP(clk), .Q(
        \input_weight[4][51] ) );
  EDFQD1 \input_weight_reg[4][50]  ( .D(data_in[50]), .E(n461), .CP(clk), .Q(
        \input_weight[4][50] ) );
  EDFQD1 \input_weight_reg[4][49]  ( .D(data_in[49]), .E(n461), .CP(clk), .Q(
        \input_weight[4][49] ) );
  EDFQD1 \input_weight_reg[4][48]  ( .D(data_in[48]), .E(n461), .CP(clk), .Q(
        \input_weight[4][48] ) );
  EDFQD1 \input_weight_reg[4][47]  ( .D(data_in[47]), .E(n461), .CP(clk), .Q(
        \input_weight[4][47] ) );
  EDFQD1 \input_weight_reg[4][46]  ( .D(data_in[46]), .E(n461), .CP(clk), .Q(
        \input_weight[4][46] ) );
  EDFQD1 \input_weight_reg[4][45]  ( .D(data_in[45]), .E(n461), .CP(clk), .Q(
        \input_weight[4][45] ) );
  EDFQD1 \input_weight_reg[4][44]  ( .D(data_in[44]), .E(n461), .CP(clk), .Q(
        \input_weight[4][44] ) );
  EDFQD1 \input_weight_reg[4][43]  ( .D(data_in[43]), .E(n461), .CP(clk), .Q(
        \input_weight[4][43] ) );
  EDFQD1 \input_weight_reg[4][42]  ( .D(data_in[42]), .E(n461), .CP(clk), .Q(
        \input_weight[4][42] ) );
  EDFQD1 \input_weight_reg[4][41]  ( .D(data_in[41]), .E(n461), .CP(clk), .Q(
        \input_weight[4][41] ) );
  EDFQD1 \input_weight_reg[4][40]  ( .D(data_in[40]), .E(n461), .CP(clk), .Q(
        \input_weight[4][40] ) );
  EDFQD1 \input_weight_reg[4][39]  ( .D(data_in[39]), .E(n461), .CP(clk), .Q(
        \input_weight[4][39] ) );
  EDFQD1 \input_weight_reg[4][38]  ( .D(data_in[38]), .E(n460), .CP(clk), .Q(
        \input_weight[4][38] ) );
  EDFQD1 \input_weight_reg[4][37]  ( .D(data_in[37]), .E(n460), .CP(clk), .Q(
        \input_weight[4][37] ) );
  EDFQD1 \input_weight_reg[4][36]  ( .D(data_in[36]), .E(n460), .CP(clk), .Q(
        \input_weight[4][36] ) );
  EDFQD1 \input_weight_reg[4][35]  ( .D(data_in[35]), .E(n460), .CP(clk), .Q(
        \input_weight[4][35] ) );
  EDFQD1 \input_weight_reg[4][34]  ( .D(data_in[34]), .E(n460), .CP(clk), .Q(
        \input_weight[4][34] ) );
  EDFQD1 \input_weight_reg[4][33]  ( .D(data_in[33]), .E(n460), .CP(clk), .Q(
        \input_weight[4][33] ) );
  EDFQD1 \input_weight_reg[4][32]  ( .D(data_in[32]), .E(n460), .CP(clk), .Q(
        \input_weight[4][32] ) );
  EDFQD1 \input_weight_reg[4][31]  ( .D(data_in[31]), .E(n460), .CP(clk), .Q(
        \input_weight[4][31] ) );
  EDFQD1 \input_weight_reg[4][30]  ( .D(data_in[30]), .E(n460), .CP(clk), .Q(
        \input_weight[4][30] ) );
  EDFQD1 \input_weight_reg[4][29]  ( .D(data_in[29]), .E(n460), .CP(clk), .Q(
        \input_weight[4][29] ) );
  EDFQD1 \input_weight_reg[4][28]  ( .D(data_in[28]), .E(n460), .CP(clk), .Q(
        \input_weight[4][28] ) );
  EDFQD1 \input_weight_reg[4][27]  ( .D(data_in[27]), .E(n460), .CP(clk), .Q(
        \input_weight[4][27] ) );
  EDFQD1 \input_weight_reg[4][26]  ( .D(data_in[26]), .E(n460), .CP(clk), .Q(
        \input_weight[4][26] ) );
  EDFQD1 \input_weight_reg[4][25]  ( .D(data_in[25]), .E(n459), .CP(clk), .Q(
        \input_weight[4][25] ) );
  EDFQD1 \input_weight_reg[4][24]  ( .D(data_in[24]), .E(n459), .CP(clk), .Q(
        \input_weight[4][24] ) );
  EDFQD1 \input_weight_reg[4][23]  ( .D(data_in[23]), .E(n459), .CP(clk), .Q(
        \input_weight[4][23] ) );
  EDFQD1 \input_weight_reg[4][22]  ( .D(data_in[22]), .E(n459), .CP(clk), .Q(
        \input_weight[4][22] ) );
  EDFQD1 \input_weight_reg[4][21]  ( .D(data_in[21]), .E(n459), .CP(clk), .Q(
        \input_weight[4][21] ) );
  EDFQD1 \input_weight_reg[4][20]  ( .D(data_in[20]), .E(n459), .CP(clk), .Q(
        \input_weight[4][20] ) );
  EDFQD1 \input_weight_reg[4][19]  ( .D(data_in[19]), .E(n459), .CP(clk), .Q(
        \input_weight[4][19] ) );
  EDFQD1 \input_weight_reg[4][18]  ( .D(data_in[18]), .E(n459), .CP(clk), .Q(
        \input_weight[4][18] ) );
  EDFQD1 \input_weight_reg[4][17]  ( .D(data_in[17]), .E(n459), .CP(clk), .Q(
        \input_weight[4][17] ) );
  EDFQD1 \input_weight_reg[4][16]  ( .D(data_in[16]), .E(n459), .CP(clk), .Q(
        \input_weight[4][16] ) );
  EDFQD1 \input_weight_reg[4][15]  ( .D(data_in[15]), .E(n459), .CP(clk), .Q(
        \input_weight[4][15] ) );
  EDFQD1 \input_weight_reg[4][14]  ( .D(data_in[14]), .E(n459), .CP(clk), .Q(
        \input_weight[4][14] ) );
  EDFQD1 \input_weight_reg[4][13]  ( .D(data_in[13]), .E(n459), .CP(clk), .Q(
        \input_weight[4][13] ) );
  EDFQD1 \input_weight_reg[4][12]  ( .D(data_in[12]), .E(n458), .CP(clk), .Q(
        \input_weight[4][12] ) );
  EDFQD1 \input_weight_reg[4][11]  ( .D(data_in[11]), .E(n458), .CP(clk), .Q(
        \input_weight[4][11] ) );
  EDFQD1 \input_weight_reg[4][10]  ( .D(data_in[10]), .E(n458), .CP(clk), .Q(
        \input_weight[4][10] ) );
  EDFQD1 \input_weight_reg[4][9]  ( .D(data_in[9]), .E(n458), .CP(clk), .Q(
        \input_weight[4][9] ) );
  EDFQD1 \input_weight_reg[4][8]  ( .D(data_in[8]), .E(n458), .CP(clk), .Q(
        \input_weight[4][8] ) );
  EDFQD1 \input_weight_reg[4][7]  ( .D(data_in[7]), .E(n458), .CP(clk), .Q(
        \input_weight[4][7] ) );
  EDFQD1 \input_weight_reg[4][6]  ( .D(data_in[6]), .E(n458), .CP(clk), .Q(
        \input_weight[4][6] ) );
  EDFQD1 \input_weight_reg[4][5]  ( .D(data_in[5]), .E(n458), .CP(clk), .Q(
        \input_weight[4][5] ) );
  EDFQD1 \input_weight_reg[4][4]  ( .D(data_in[4]), .E(n458), .CP(clk), .Q(
        \input_weight[4][4] ) );
  EDFQD1 \input_weight_reg[4][3]  ( .D(data_in[3]), .E(n458), .CP(clk), .Q(
        \input_weight[4][3] ) );
  EDFQD1 \input_weight_reg[4][2]  ( .D(data_in[2]), .E(n458), .CP(clk), .Q(
        \input_weight[4][2] ) );
  EDFQD1 \input_weight_reg[4][1]  ( .D(data_in[1]), .E(n458), .CP(clk), .Q(
        \input_weight[4][1] ) );
  EDFQD1 \input_weight_reg[4][0]  ( .D(data_in[0]), .E(n458), .CP(clk), .Q(
        \input_weight[4][0] ) );
  EDFQD1 \input_bias_reg[3][5]  ( .D(data_in[5]), .E(N480), .CP(clk), .Q(
        \input_bias[3][5] ) );
  EDFQD1 \input_bias_reg[3][4]  ( .D(data_in[4]), .E(N480), .CP(clk), .Q(
        \input_bias[3][4] ) );
  EDFQD1 \input_bias_reg[3][3]  ( .D(data_in[3]), .E(N480), .CP(clk), .Q(
        \input_bias[3][3] ) );
  EDFQD1 \input_bias_reg[3][2]  ( .D(data_in[2]), .E(N480), .CP(clk), .Q(
        \input_bias[3][2] ) );
  EDFQD1 \input_bias_reg[3][1]  ( .D(data_in[1]), .E(N480), .CP(clk), .Q(
        \input_bias[3][1] ) );
  EDFQD1 \input_bias_reg[3][0]  ( .D(data_in[0]), .E(N480), .CP(clk), .Q(
        \input_bias[3][0] ) );
  EDFQD1 \input_bias_reg[1][5]  ( .D(data_in[5]), .E(N478), .CP(clk), .Q(
        \input_bias[1][5] ) );
  EDFQD1 \input_bias_reg[1][4]  ( .D(data_in[4]), .E(N478), .CP(clk), .Q(
        \input_bias[1][4] ) );
  EDFQD1 \input_bias_reg[1][3]  ( .D(data_in[3]), .E(N478), .CP(clk), .Q(
        \input_bias[1][3] ) );
  EDFQD1 \input_bias_reg[1][2]  ( .D(data_in[2]), .E(N478), .CP(clk), .Q(
        \input_bias[1][2] ) );
  EDFQD1 \input_bias_reg[1][1]  ( .D(data_in[1]), .E(N478), .CP(clk), .Q(
        \input_bias[1][1] ) );
  EDFQD1 \input_bias_reg[1][0]  ( .D(data_in[0]), .E(N478), .CP(clk), .Q(
        \input_bias[1][0] ) );
  EDFQD1 \input_bias_reg[6][5]  ( .D(data_in[5]), .E(N483), .CP(clk), .Q(
        \input_bias[6][5] ) );
  EDFQD1 \input_bias_reg[6][4]  ( .D(data_in[4]), .E(N483), .CP(clk), .Q(
        \input_bias[6][4] ) );
  EDFQD1 \input_bias_reg[6][3]  ( .D(data_in[3]), .E(N483), .CP(clk), .Q(
        \input_bias[6][3] ) );
  EDFQD1 \input_bias_reg[6][2]  ( .D(data_in[2]), .E(N483), .CP(clk), .Q(
        \input_bias[6][2] ) );
  EDFQD1 \input_bias_reg[6][1]  ( .D(data_in[1]), .E(N483), .CP(clk), .Q(
        \input_bias[6][1] ) );
  EDFQD1 \input_bias_reg[6][0]  ( .D(data_in[0]), .E(N483), .CP(clk), .Q(
        \input_bias[6][0] ) );
  EDFQD1 \input_bias_reg[4][5]  ( .D(data_in[5]), .E(N481), .CP(clk), .Q(
        \input_bias[4][5] ) );
  EDFQD1 \input_bias_reg[4][4]  ( .D(data_in[4]), .E(N481), .CP(clk), .Q(
        \input_bias[4][4] ) );
  EDFQD1 \input_bias_reg[4][3]  ( .D(data_in[3]), .E(N481), .CP(clk), .Q(
        \input_bias[4][3] ) );
  EDFQD1 \input_bias_reg[4][2]  ( .D(data_in[2]), .E(N481), .CP(clk), .Q(
        \input_bias[4][2] ) );
  EDFQD1 \input_bias_reg[4][1]  ( .D(data_in[1]), .E(N481), .CP(clk), .Q(
        \input_bias[4][1] ) );
  EDFQD1 \input_bias_reg[4][0]  ( .D(data_in[0]), .E(N481), .CP(clk), .Q(
        \input_bias[4][0] ) );
  EDFQD1 \input_bias_reg[0][5]  ( .D(data_in[5]), .E(N477), .CP(clk), .Q(
        \input_bias[0][5] ) );
  EDFQD1 \input_bias_reg[0][4]  ( .D(data_in[4]), .E(N477), .CP(clk), .Q(
        \input_bias[0][4] ) );
  EDFQD1 \input_bias_reg[0][3]  ( .D(data_in[3]), .E(N477), .CP(clk), .Q(
        \input_bias[0][3] ) );
  EDFQD1 \input_bias_reg[0][2]  ( .D(data_in[2]), .E(N477), .CP(clk), .Q(
        \input_bias[0][2] ) );
  EDFQD1 \input_bias_reg[0][1]  ( .D(data_in[1]), .E(N477), .CP(clk), .Q(
        \input_bias[0][1] ) );
  EDFQD1 \input_bias_reg[0][0]  ( .D(data_in[0]), .E(N477), .CP(clk), .Q(
        \input_bias[0][0] ) );
  EDFQD1 \input_bias_reg[2][5]  ( .D(data_in[5]), .E(N479), .CP(clk), .Q(
        \input_bias[2][5] ) );
  EDFQD1 \input_bias_reg[2][4]  ( .D(data_in[4]), .E(N479), .CP(clk), .Q(
        \input_bias[2][4] ) );
  EDFQD1 \input_bias_reg[2][3]  ( .D(data_in[3]), .E(N479), .CP(clk), .Q(
        \input_bias[2][3] ) );
  EDFQD1 \input_bias_reg[2][2]  ( .D(data_in[2]), .E(N479), .CP(clk), .Q(
        \input_bias[2][2] ) );
  EDFQD1 \input_bias_reg[2][1]  ( .D(data_in[1]), .E(N479), .CP(clk), .Q(
        \input_bias[2][1] ) );
  EDFQD1 \input_bias_reg[2][0]  ( .D(data_in[0]), .E(N479), .CP(clk), .Q(
        \input_bias[2][0] ) );
  EDFQD1 \input_bias_reg[5][5]  ( .D(data_in[5]), .E(N482), .CP(clk), .Q(
        \input_bias[5][5] ) );
  EDFQD1 \input_bias_reg[5][4]  ( .D(data_in[4]), .E(N482), .CP(clk), .Q(
        \input_bias[5][4] ) );
  EDFQD1 \input_bias_reg[5][3]  ( .D(data_in[3]), .E(N482), .CP(clk), .Q(
        \input_bias[5][3] ) );
  EDFQD1 \input_bias_reg[5][2]  ( .D(data_in[2]), .E(N482), .CP(clk), .Q(
        \input_bias[5][2] ) );
  EDFQD1 \input_bias_reg[5][1]  ( .D(data_in[1]), .E(N482), .CP(clk), .Q(
        \input_bias[5][1] ) );
  EDFQD1 \input_bias_reg[5][0]  ( .D(data_in[0]), .E(N482), .CP(clk), .Q(
        \input_bias[5][0] ) );
  EDFQD1 \input_bias_reg[7][5]  ( .D(data_in[5]), .E(N484), .CP(clk), .Q(
        \input_bias[7][5] ) );
  EDFQD1 \input_bias_reg[7][4]  ( .D(data_in[4]), .E(N484), .CP(clk), .Q(
        \input_bias[7][4] ) );
  EDFQD1 \input_bias_reg[7][3]  ( .D(data_in[3]), .E(N484), .CP(clk), .Q(
        \input_bias[7][3] ) );
  EDFQD1 \input_bias_reg[7][2]  ( .D(data_in[2]), .E(N484), .CP(clk), .Q(
        \input_bias[7][2] ) );
  EDFQD1 \input_bias_reg[7][1]  ( .D(data_in[1]), .E(N484), .CP(clk), .Q(
        \input_bias[7][1] ) );
  EDFQD1 \input_bias_reg[7][0]  ( .D(data_in[0]), .E(N484), .CP(clk), .Q(
        \input_bias[7][0] ) );
  EDFQD1 \mem_nxt_state_reg[3]  ( .D(N317), .E(N312), .CP(clk), .Q(
        mem_nxt_state[3]) );
  EDFQD1 \mem_nxt_state_reg[1]  ( .D(N315), .E(N312), .CP(clk), .Q(
        mem_nxt_state[1]) );
  EDFQD1 \input_bias_reg[6][15]  ( .D(data_in[15]), .E(N483), .CP(clk), .Q(
        \input_bias[6][15] ) );
  EDFQD1 \input_bias_reg[6][14]  ( .D(data_in[14]), .E(N483), .CP(clk), .Q(
        \input_bias[6][14] ) );
  EDFQD1 \input_bias_reg[6][13]  ( .D(data_in[13]), .E(N483), .CP(clk), .Q(
        \input_bias[6][13] ) );
  EDFQD1 \input_bias_reg[6][12]  ( .D(data_in[12]), .E(N483), .CP(clk), .Q(
        \input_bias[6][12] ) );
  EDFQD1 \input_bias_reg[6][11]  ( .D(data_in[11]), .E(N483), .CP(clk), .Q(
        \input_bias[6][11] ) );
  EDFQD1 \input_bias_reg[6][10]  ( .D(data_in[10]), .E(N483), .CP(clk), .Q(
        \input_bias[6][10] ) );
  EDFQD1 \input_bias_reg[6][9]  ( .D(data_in[9]), .E(N483), .CP(clk), .Q(
        \input_bias[6][9] ) );
  EDFQD1 \input_bias_reg[6][8]  ( .D(data_in[8]), .E(N483), .CP(clk), .Q(
        \input_bias[6][8] ) );
  EDFQD1 \input_bias_reg[6][7]  ( .D(data_in[7]), .E(N483), .CP(clk), .Q(
        \input_bias[6][7] ) );
  EDFQD1 \input_bias_reg[6][6]  ( .D(data_in[6]), .E(N483), .CP(clk), .Q(
        \input_bias[6][6] ) );
  EDFQD1 \mem_nxt_state_reg[2]  ( .D(\U3/U1/Z_5 ), .E(N312), .CP(clk), .Q(
        mem_nxt_state[2]) );
  EDFQD1 \mem_nxt_state_reg[0]  ( .D(N314), .E(N312), .CP(clk), .Q(
        mem_nxt_state[0]) );
  EDFQD1 \input_bias_reg[2][15]  ( .D(data_in[15]), .E(N479), .CP(clk), .Q(
        \input_bias[2][15] ) );
  EDFQD1 \input_bias_reg[2][14]  ( .D(data_in[14]), .E(N479), .CP(clk), .Q(
        \input_bias[2][14] ) );
  EDFQD1 \input_bias_reg[2][13]  ( .D(data_in[13]), .E(N479), .CP(clk), .Q(
        \input_bias[2][13] ) );
  EDFQD1 \input_bias_reg[2][12]  ( .D(data_in[12]), .E(N479), .CP(clk), .Q(
        \input_bias[2][12] ) );
  EDFQD1 \input_bias_reg[2][11]  ( .D(data_in[11]), .E(N479), .CP(clk), .Q(
        \input_bias[2][11] ) );
  EDFQD1 \input_bias_reg[2][10]  ( .D(data_in[10]), .E(N479), .CP(clk), .Q(
        \input_bias[2][10] ) );
  EDFQD1 \input_bias_reg[2][9]  ( .D(data_in[9]), .E(N479), .CP(clk), .Q(
        \input_bias[2][9] ) );
  EDFQD1 \input_bias_reg[2][8]  ( .D(data_in[8]), .E(N479), .CP(clk), .Q(
        \input_bias[2][8] ) );
  EDFQD1 \input_bias_reg[2][7]  ( .D(data_in[7]), .E(N479), .CP(clk), .Q(
        \input_bias[2][7] ) );
  EDFQD1 \input_bias_reg[2][6]  ( .D(data_in[6]), .E(N479), .CP(clk), .Q(
        \input_bias[2][6] ) );
  EDFQD1 \input_bias_reg[4][15]  ( .D(data_in[15]), .E(N481), .CP(clk), .Q(
        \input_bias[4][15] ) );
  EDFQD1 \input_bias_reg[4][14]  ( .D(data_in[14]), .E(N481), .CP(clk), .Q(
        \input_bias[4][14] ) );
  EDFQD1 \input_bias_reg[4][13]  ( .D(data_in[13]), .E(N481), .CP(clk), .Q(
        \input_bias[4][13] ) );
  EDFQD1 \input_bias_reg[4][12]  ( .D(data_in[12]), .E(N481), .CP(clk), .Q(
        \input_bias[4][12] ) );
  EDFQD1 \input_bias_reg[4][11]  ( .D(data_in[11]), .E(N481), .CP(clk), .Q(
        \input_bias[4][11] ) );
  EDFQD1 \input_bias_reg[4][10]  ( .D(data_in[10]), .E(N481), .CP(clk), .Q(
        \input_bias[4][10] ) );
  EDFQD1 \input_bias_reg[4][9]  ( .D(data_in[9]), .E(N481), .CP(clk), .Q(
        \input_bias[4][9] ) );
  EDFQD1 \input_bias_reg[4][8]  ( .D(data_in[8]), .E(N481), .CP(clk), .Q(
        \input_bias[4][8] ) );
  EDFQD1 \input_bias_reg[4][7]  ( .D(data_in[7]), .E(N481), .CP(clk), .Q(
        \input_bias[4][7] ) );
  EDFQD1 \input_bias_reg[4][6]  ( .D(data_in[6]), .E(N481), .CP(clk), .Q(
        \input_bias[4][6] ) );
  EDFQD1 \input_bias_reg[0][15]  ( .D(data_in[15]), .E(N477), .CP(clk), .Q(
        \input_bias[0][15] ) );
  EDFQD1 \input_bias_reg[0][14]  ( .D(data_in[14]), .E(N477), .CP(clk), .Q(
        \input_bias[0][14] ) );
  EDFQD1 \input_bias_reg[0][13]  ( .D(data_in[13]), .E(N477), .CP(clk), .Q(
        \input_bias[0][13] ) );
  EDFQD1 \input_bias_reg[0][12]  ( .D(data_in[12]), .E(N477), .CP(clk), .Q(
        \input_bias[0][12] ) );
  EDFQD1 \input_bias_reg[0][11]  ( .D(data_in[11]), .E(N477), .CP(clk), .Q(
        \input_bias[0][11] ) );
  EDFQD1 \input_bias_reg[0][10]  ( .D(data_in[10]), .E(N477), .CP(clk), .Q(
        \input_bias[0][10] ) );
  EDFQD1 \input_bias_reg[0][9]  ( .D(data_in[9]), .E(N477), .CP(clk), .Q(
        \input_bias[0][9] ) );
  EDFQD1 \input_bias_reg[0][8]  ( .D(data_in[8]), .E(N477), .CP(clk), .Q(
        \input_bias[0][8] ) );
  EDFQD1 \input_bias_reg[0][7]  ( .D(data_in[7]), .E(N477), .CP(clk), .Q(
        \input_bias[0][7] ) );
  EDFQD1 \input_bias_reg[0][6]  ( .D(data_in[6]), .E(N477), .CP(clk), .Q(
        \input_bias[0][6] ) );
  EDFQD1 \input_bias_reg[7][15]  ( .D(data_in[15]), .E(N484), .CP(clk), .Q(
        \input_bias[7][15] ) );
  EDFQD1 \input_bias_reg[7][14]  ( .D(data_in[14]), .E(N484), .CP(clk), .Q(
        \input_bias[7][14] ) );
  EDFQD1 \input_bias_reg[7][13]  ( .D(data_in[13]), .E(N484), .CP(clk), .Q(
        \input_bias[7][13] ) );
  EDFQD1 \input_bias_reg[7][12]  ( .D(data_in[12]), .E(N484), .CP(clk), .Q(
        \input_bias[7][12] ) );
  EDFQD1 \input_bias_reg[7][11]  ( .D(data_in[11]), .E(N484), .CP(clk), .Q(
        \input_bias[7][11] ) );
  EDFQD1 \input_bias_reg[7][10]  ( .D(data_in[10]), .E(N484), .CP(clk), .Q(
        \input_bias[7][10] ) );
  EDFQD1 \input_bias_reg[7][9]  ( .D(data_in[9]), .E(N484), .CP(clk), .Q(
        \input_bias[7][9] ) );
  EDFQD1 \input_bias_reg[7][8]  ( .D(data_in[8]), .E(N484), .CP(clk), .Q(
        \input_bias[7][8] ) );
  EDFQD1 \input_bias_reg[7][7]  ( .D(data_in[7]), .E(N484), .CP(clk), .Q(
        \input_bias[7][7] ) );
  EDFQD1 \input_bias_reg[7][6]  ( .D(data_in[6]), .E(N484), .CP(clk), .Q(
        \input_bias[7][6] ) );
  EDFQD1 \input_bias_reg[5][15]  ( .D(data_in[15]), .E(N482), .CP(clk), .Q(
        \input_bias[5][15] ) );
  EDFQD1 \input_bias_reg[5][14]  ( .D(data_in[14]), .E(N482), .CP(clk), .Q(
        \input_bias[5][14] ) );
  EDFQD1 \input_bias_reg[5][13]  ( .D(data_in[13]), .E(N482), .CP(clk), .Q(
        \input_bias[5][13] ) );
  EDFQD1 \input_bias_reg[5][12]  ( .D(data_in[12]), .E(N482), .CP(clk), .Q(
        \input_bias[5][12] ) );
  EDFQD1 \input_bias_reg[5][11]  ( .D(data_in[11]), .E(N482), .CP(clk), .Q(
        \input_bias[5][11] ) );
  EDFQD1 \input_bias_reg[5][10]  ( .D(data_in[10]), .E(N482), .CP(clk), .Q(
        \input_bias[5][10] ) );
  EDFQD1 \input_bias_reg[5][9]  ( .D(data_in[9]), .E(N482), .CP(clk), .Q(
        \input_bias[5][9] ) );
  EDFQD1 \input_bias_reg[5][8]  ( .D(data_in[8]), .E(N482), .CP(clk), .Q(
        \input_bias[5][8] ) );
  EDFQD1 \input_bias_reg[5][7]  ( .D(data_in[7]), .E(N482), .CP(clk), .Q(
        \input_bias[5][7] ) );
  EDFQD1 \input_bias_reg[5][6]  ( .D(data_in[6]), .E(N482), .CP(clk), .Q(
        \input_bias[5][6] ) );
  EDFQD1 \input_bias_reg[1][15]  ( .D(data_in[15]), .E(N478), .CP(clk), .Q(
        \input_bias[1][15] ) );
  EDFQD1 \input_bias_reg[1][14]  ( .D(data_in[14]), .E(N478), .CP(clk), .Q(
        \input_bias[1][14] ) );
  EDFQD1 \input_bias_reg[1][13]  ( .D(data_in[13]), .E(N478), .CP(clk), .Q(
        \input_bias[1][13] ) );
  EDFQD1 \input_bias_reg[1][12]  ( .D(data_in[12]), .E(N478), .CP(clk), .Q(
        \input_bias[1][12] ) );
  EDFQD1 \input_bias_reg[1][11]  ( .D(data_in[11]), .E(N478), .CP(clk), .Q(
        \input_bias[1][11] ) );
  EDFQD1 \input_bias_reg[1][10]  ( .D(data_in[10]), .E(N478), .CP(clk), .Q(
        \input_bias[1][10] ) );
  EDFQD1 \input_bias_reg[1][9]  ( .D(data_in[9]), .E(N478), .CP(clk), .Q(
        \input_bias[1][9] ) );
  EDFQD1 \input_bias_reg[1][8]  ( .D(data_in[8]), .E(N478), .CP(clk), .Q(
        \input_bias[1][8] ) );
  EDFQD1 \input_bias_reg[1][7]  ( .D(data_in[7]), .E(N478), .CP(clk), .Q(
        \input_bias[1][7] ) );
  EDFQD1 \input_bias_reg[1][6]  ( .D(data_in[6]), .E(N478), .CP(clk), .Q(
        \input_bias[1][6] ) );
  EDFQD1 \input_bias_reg[3][15]  ( .D(data_in[15]), .E(N480), .CP(clk), .Q(
        \input_bias[3][15] ) );
  EDFQD1 \input_bias_reg[3][14]  ( .D(data_in[14]), .E(N480), .CP(clk), .Q(
        \input_bias[3][14] ) );
  EDFQD1 \input_bias_reg[3][13]  ( .D(data_in[13]), .E(N480), .CP(clk), .Q(
        \input_bias[3][13] ) );
  EDFQD1 \input_bias_reg[3][12]  ( .D(data_in[12]), .E(N480), .CP(clk), .Q(
        \input_bias[3][12] ) );
  EDFQD1 \input_bias_reg[3][11]  ( .D(data_in[11]), .E(N480), .CP(clk), .Q(
        \input_bias[3][11] ) );
  EDFQD1 \input_bias_reg[3][10]  ( .D(data_in[10]), .E(N480), .CP(clk), .Q(
        \input_bias[3][10] ) );
  EDFQD1 \input_bias_reg[3][9]  ( .D(data_in[9]), .E(N480), .CP(clk), .Q(
        \input_bias[3][9] ) );
  EDFQD1 \input_bias_reg[3][8]  ( .D(data_in[8]), .E(N480), .CP(clk), .Q(
        \input_bias[3][8] ) );
  EDFQD1 \input_bias_reg[3][7]  ( .D(data_in[7]), .E(N480), .CP(clk), .Q(
        \input_bias[3][7] ) );
  EDFQD1 \input_bias_reg[3][6]  ( .D(data_in[6]), .E(N480), .CP(clk), .Q(
        \input_bias[3][6] ) );
  NR2XD0 U309 ( .A1(n537), .A2(n538), .ZN(N484) );
  NR2XD0 U310 ( .A1(n537), .A2(n540), .ZN(N482) );
  NR2XD0 U311 ( .A1(n537), .A2(n543), .ZN(N479) );
  NR2XD0 U312 ( .A1(n537), .A2(n544), .ZN(N477) );
  NR2XD0 U313 ( .A1(n537), .A2(n541), .ZN(N481) );
  NR2XD0 U314 ( .A1(n537), .A2(n539), .ZN(N483) );
  NR2XD0 U315 ( .A1(n537), .A2(n536), .ZN(N478) );
  NR2XD0 U316 ( .A1(n537), .A2(n542), .ZN(N480) );
  ND4D2 U317 ( .A1(n564), .A2(n546), .A3(n568), .A4(n535), .ZN(N312) );
  CKBD1 U318 ( .I(n472), .Z(n458) );
  CKBD1 U319 ( .I(n472), .Z(n459) );
  CKBD1 U320 ( .I(n471), .Z(n460) );
  CKBD1 U321 ( .I(n471), .Z(n461) );
  CKBD1 U322 ( .I(n470), .Z(n462) );
  CKBD1 U323 ( .I(n470), .Z(n463) );
  CKBD1 U324 ( .I(n469), .Z(n464) );
  CKBD1 U325 ( .I(n469), .Z(n465) );
  CKBD1 U326 ( .I(n468), .Z(n466) );
  CKBD1 U327 ( .I(n352), .Z(n338) );
  CKBD1 U328 ( .I(n352), .Z(n339) );
  CKBD1 U329 ( .I(n351), .Z(n340) );
  CKBD1 U330 ( .I(n351), .Z(n341) );
  CKBD1 U331 ( .I(n350), .Z(n342) );
  CKBD1 U332 ( .I(n350), .Z(n343) );
  CKBD1 U333 ( .I(n349), .Z(n344) );
  CKBD1 U334 ( .I(n349), .Z(n345) );
  CKBD1 U335 ( .I(n348), .Z(n346) );
  CKBD1 U336 ( .I(n468), .Z(n467) );
  CKBD1 U337 ( .I(n348), .Z(n347) );
  CKBD1 U338 ( .I(N438), .Z(n472) );
  CKBD1 U339 ( .I(N438), .Z(n471) );
  CKBD1 U340 ( .I(N438), .Z(n470) );
  CKBD1 U341 ( .I(N438), .Z(n469) );
  CKBD1 U342 ( .I(N438), .Z(n468) );
  CKBD1 U343 ( .I(N454), .Z(n352) );
  CKBD1 U344 ( .I(N454), .Z(n351) );
  CKBD1 U345 ( .I(N454), .Z(n350) );
  CKBD1 U346 ( .I(N454), .Z(n349) );
  CKBD1 U347 ( .I(N454), .Z(n348) );
  CKBD1 U348 ( .I(n487), .Z(n473) );
  CKBD1 U349 ( .I(n487), .Z(n474) );
  CKBD1 U350 ( .I(n486), .Z(n475) );
  CKBD1 U351 ( .I(n486), .Z(n476) );
  CKBD1 U352 ( .I(n485), .Z(n477) );
  CKBD1 U353 ( .I(n485), .Z(n478) );
  CKBD1 U354 ( .I(n484), .Z(n479) );
  CKBD1 U355 ( .I(n484), .Z(n480) );
  CKBD1 U356 ( .I(n483), .Z(n481) );
  CKBD1 U357 ( .I(n367), .Z(n353) );
  CKBD1 U358 ( .I(n367), .Z(n354) );
  CKBD1 U359 ( .I(n366), .Z(n355) );
  CKBD1 U360 ( .I(n366), .Z(n356) );
  CKBD1 U361 ( .I(n365), .Z(n357) );
  CKBD1 U362 ( .I(n365), .Z(n358) );
  CKBD1 U363 ( .I(n364), .Z(n359) );
  CKBD1 U364 ( .I(n364), .Z(n360) );
  CKBD1 U365 ( .I(n363), .Z(n361) );
  CKBD1 U366 ( .I(n517), .Z(n503) );
  CKBD1 U367 ( .I(n517), .Z(n504) );
  CKBD1 U368 ( .I(n516), .Z(n505) );
  CKBD1 U369 ( .I(n516), .Z(n506) );
  CKBD1 U370 ( .I(n515), .Z(n507) );
  CKBD1 U371 ( .I(n515), .Z(n508) );
  CKBD1 U372 ( .I(n514), .Z(n509) );
  CKBD1 U373 ( .I(n514), .Z(n510) );
  CKBD1 U374 ( .I(n513), .Z(n511) );
  CKBD1 U375 ( .I(n397), .Z(n383) );
  CKBD1 U376 ( .I(n397), .Z(n384) );
  CKBD1 U377 ( .I(n396), .Z(n385) );
  CKBD1 U378 ( .I(n396), .Z(n386) );
  CKBD1 U379 ( .I(n395), .Z(n387) );
  CKBD1 U380 ( .I(n395), .Z(n388) );
  CKBD1 U381 ( .I(n394), .Z(n389) );
  CKBD1 U382 ( .I(n394), .Z(n390) );
  CKBD1 U383 ( .I(n393), .Z(n391) );
  CKBD1 U384 ( .I(n457), .Z(n443) );
  CKBD1 U385 ( .I(n457), .Z(n444) );
  CKBD1 U386 ( .I(n456), .Z(n445) );
  CKBD1 U387 ( .I(n456), .Z(n446) );
  CKBD1 U388 ( .I(n455), .Z(n447) );
  CKBD1 U389 ( .I(n455), .Z(n448) );
  CKBD1 U390 ( .I(n454), .Z(n449) );
  CKBD1 U391 ( .I(n454), .Z(n450) );
  CKBD1 U392 ( .I(n453), .Z(n451) );
  CKBD1 U393 ( .I(n337), .Z(n323) );
  CKBD1 U394 ( .I(n337), .Z(n324) );
  CKBD1 U395 ( .I(n336), .Z(n325) );
  CKBD1 U396 ( .I(n336), .Z(n326) );
  CKBD1 U397 ( .I(n335), .Z(n327) );
  CKBD1 U398 ( .I(n335), .Z(n328) );
  CKBD1 U399 ( .I(n334), .Z(n329) );
  CKBD1 U400 ( .I(n334), .Z(n330) );
  CKBD1 U401 ( .I(n333), .Z(n331) );
  CKBD1 U402 ( .I(n427), .Z(n413) );
  CKBD1 U403 ( .I(n427), .Z(n414) );
  CKBD1 U404 ( .I(n426), .Z(n415) );
  CKBD1 U405 ( .I(n426), .Z(n416) );
  CKBD1 U406 ( .I(n425), .Z(n417) );
  CKBD1 U407 ( .I(n425), .Z(n418) );
  CKBD1 U408 ( .I(n424), .Z(n419) );
  CKBD1 U409 ( .I(n424), .Z(n420) );
  CKBD1 U410 ( .I(n423), .Z(n421) );
  CKBD1 U411 ( .I(n307), .Z(n293) );
  CKBD1 U412 ( .I(n307), .Z(n294) );
  CKBD1 U413 ( .I(n306), .Z(n295) );
  CKBD1 U414 ( .I(n306), .Z(n296) );
  CKBD1 U415 ( .I(n305), .Z(n297) );
  CKBD1 U416 ( .I(n305), .Z(n298) );
  CKBD1 U417 ( .I(n304), .Z(n299) );
  CKBD1 U418 ( .I(n304), .Z(n300) );
  CKBD1 U419 ( .I(n303), .Z(n301) );
  CKBD1 U420 ( .I(n532), .Z(n518) );
  CKBD1 U421 ( .I(n532), .Z(n519) );
  CKBD1 U422 ( .I(n531), .Z(n520) );
  CKBD1 U423 ( .I(n531), .Z(n521) );
  CKBD1 U424 ( .I(n530), .Z(n522) );
  CKBD1 U425 ( .I(n530), .Z(n523) );
  CKBD1 U426 ( .I(n529), .Z(n524) );
  CKBD1 U427 ( .I(n529), .Z(n525) );
  CKBD1 U428 ( .I(n528), .Z(n526) );
  CKBD1 U429 ( .I(n412), .Z(n398) );
  CKBD1 U430 ( .I(n412), .Z(n399) );
  CKBD1 U431 ( .I(n411), .Z(n400) );
  CKBD1 U432 ( .I(n411), .Z(n401) );
  CKBD1 U433 ( .I(n410), .Z(n402) );
  CKBD1 U434 ( .I(n410), .Z(n403) );
  CKBD1 U435 ( .I(n409), .Z(n404) );
  CKBD1 U436 ( .I(n409), .Z(n405) );
  CKBD1 U437 ( .I(n408), .Z(n406) );
  CKBD1 U438 ( .I(n502), .Z(n488) );
  CKBD1 U439 ( .I(n502), .Z(n489) );
  CKBD1 U440 ( .I(n501), .Z(n490) );
  CKBD1 U441 ( .I(n501), .Z(n491) );
  CKBD1 U442 ( .I(n500), .Z(n492) );
  CKBD1 U443 ( .I(n500), .Z(n493) );
  CKBD1 U444 ( .I(n499), .Z(n494) );
  CKBD1 U445 ( .I(n499), .Z(n495) );
  CKBD1 U446 ( .I(n498), .Z(n496) );
  CKBD1 U447 ( .I(n382), .Z(n368) );
  CKBD1 U448 ( .I(n382), .Z(n369) );
  CKBD1 U449 ( .I(n381), .Z(n370) );
  CKBD1 U450 ( .I(n381), .Z(n371) );
  CKBD1 U451 ( .I(n380), .Z(n372) );
  CKBD1 U452 ( .I(n380), .Z(n373) );
  CKBD1 U453 ( .I(n379), .Z(n374) );
  CKBD1 U454 ( .I(n379), .Z(n375) );
  CKBD1 U455 ( .I(n378), .Z(n376) );
  CKBD1 U456 ( .I(n277), .Z(n264) );
  CKBD1 U457 ( .I(n277), .Z(n263) );
  CKBD1 U458 ( .I(n292), .Z(n279) );
  CKBD1 U459 ( .I(n292), .Z(n278) );
  CKBD1 U460 ( .I(n322), .Z(n308) );
  CKBD1 U461 ( .I(n322), .Z(n309) );
  CKBD1 U462 ( .I(n321), .Z(n310) );
  CKBD1 U463 ( .I(n321), .Z(n311) );
  CKBD1 U464 ( .I(n320), .Z(n312) );
  CKBD1 U465 ( .I(n320), .Z(n313) );
  CKBD1 U466 ( .I(n319), .Z(n314) );
  CKBD1 U467 ( .I(n319), .Z(n315) );
  CKBD1 U468 ( .I(n318), .Z(n316) );
  CKBD1 U469 ( .I(n442), .Z(n428) );
  CKBD1 U470 ( .I(n442), .Z(n429) );
  CKBD1 U471 ( .I(n441), .Z(n430) );
  CKBD1 U472 ( .I(n441), .Z(n431) );
  CKBD1 U473 ( .I(n440), .Z(n432) );
  CKBD1 U474 ( .I(n440), .Z(n433) );
  CKBD1 U475 ( .I(n439), .Z(n434) );
  CKBD1 U476 ( .I(n439), .Z(n435) );
  CKBD1 U477 ( .I(n438), .Z(n436) );
  CKBD1 U478 ( .I(n276), .Z(n265) );
  CKBD1 U479 ( .I(n276), .Z(n266) );
  CKBD1 U480 ( .I(n275), .Z(n267) );
  CKBD1 U481 ( .I(n275), .Z(n268) );
  CKBD1 U482 ( .I(n274), .Z(n269) );
  CKBD1 U483 ( .I(n274), .Z(n270) );
  CKBD1 U484 ( .I(n273), .Z(n271) );
  CKBD1 U485 ( .I(n291), .Z(n280) );
  CKBD1 U486 ( .I(n291), .Z(n281) );
  CKBD1 U487 ( .I(n290), .Z(n282) );
  CKBD1 U488 ( .I(n290), .Z(n283) );
  CKBD1 U489 ( .I(n289), .Z(n284) );
  CKBD1 U490 ( .I(n289), .Z(n285) );
  CKBD1 U491 ( .I(n288), .Z(n286) );
  CKBD1 U492 ( .I(n483), .Z(n482) );
  CKBD1 U493 ( .I(n363), .Z(n362) );
  CKBD1 U494 ( .I(n513), .Z(n512) );
  CKBD1 U495 ( .I(n393), .Z(n392) );
  CKBD1 U496 ( .I(n453), .Z(n452) );
  CKBD1 U497 ( .I(n333), .Z(n332) );
  CKBD1 U498 ( .I(n423), .Z(n422) );
  CKBD1 U499 ( .I(n303), .Z(n302) );
  CKBD1 U500 ( .I(n528), .Z(n527) );
  CKBD1 U501 ( .I(n408), .Z(n407) );
  CKBD1 U502 ( .I(n498), .Z(n497) );
  CKBD1 U503 ( .I(n378), .Z(n377) );
  CKBD1 U504 ( .I(n318), .Z(n317) );
  CKBD1 U505 ( .I(n438), .Z(n437) );
  CKBD1 U506 ( .I(n273), .Z(n272) );
  CKBD1 U507 ( .I(n288), .Z(n287) );
  CKBD1 U508 ( .I(N440), .Z(n457) );
  CKBD1 U509 ( .I(N440), .Z(n456) );
  CKBD1 U510 ( .I(N440), .Z(n455) );
  CKBD1 U511 ( .I(N440), .Z(n454) );
  CKBD1 U512 ( .I(N440), .Z(n453) );
  CKBD1 U513 ( .I(N456), .Z(n337) );
  CKBD1 U514 ( .I(N456), .Z(n336) );
  CKBD1 U515 ( .I(N456), .Z(n335) );
  CKBD1 U516 ( .I(N456), .Z(n334) );
  CKBD1 U517 ( .I(N456), .Z(n333) );
  CKBD1 U518 ( .I(N430), .Z(n532) );
  CKBD1 U519 ( .I(N430), .Z(n531) );
  CKBD1 U520 ( .I(N430), .Z(n530) );
  CKBD1 U521 ( .I(N430), .Z(n529) );
  CKBD1 U522 ( .I(N430), .Z(n528) );
  CKBD1 U523 ( .I(N446), .Z(n412) );
  CKBD1 U524 ( .I(N446), .Z(n411) );
  CKBD1 U525 ( .I(N446), .Z(n410) );
  CKBD1 U526 ( .I(N446), .Z(n409) );
  CKBD1 U527 ( .I(N446), .Z(n408) );
  CKBD1 U528 ( .I(N458), .Z(n322) );
  CKBD1 U529 ( .I(N458), .Z(n321) );
  CKBD1 U530 ( .I(N458), .Z(n320) );
  CKBD1 U531 ( .I(N458), .Z(n319) );
  CKBD1 U532 ( .I(N458), .Z(n318) );
  CKBD1 U533 ( .I(N442), .Z(n442) );
  CKBD1 U534 ( .I(N442), .Z(n441) );
  CKBD1 U535 ( .I(N442), .Z(n440) );
  CKBD1 U536 ( .I(N442), .Z(n439) );
  CKBD1 U537 ( .I(N442), .Z(n438) );
  CKBD1 U538 ( .I(N436), .Z(n487) );
  CKBD1 U539 ( .I(N436), .Z(n486) );
  CKBD1 U540 ( .I(N436), .Z(n485) );
  CKBD1 U541 ( .I(N436), .Z(n484) );
  CKBD1 U542 ( .I(N436), .Z(n483) );
  CKBD1 U543 ( .I(N452), .Z(n367) );
  CKBD1 U544 ( .I(N452), .Z(n366) );
  CKBD1 U545 ( .I(N452), .Z(n365) );
  CKBD1 U546 ( .I(N452), .Z(n364) );
  CKBD1 U547 ( .I(N452), .Z(n363) );
  CKBD1 U548 ( .I(N432), .Z(n517) );
  CKBD1 U549 ( .I(N432), .Z(n516) );
  CKBD1 U550 ( .I(N432), .Z(n515) );
  CKBD1 U551 ( .I(N432), .Z(n514) );
  CKBD1 U552 ( .I(N432), .Z(n513) );
  CKBD1 U553 ( .I(N448), .Z(n397) );
  CKBD1 U554 ( .I(N448), .Z(n396) );
  CKBD1 U555 ( .I(N448), .Z(n395) );
  CKBD1 U556 ( .I(N448), .Z(n394) );
  CKBD1 U557 ( .I(N448), .Z(n393) );
  CKBD1 U558 ( .I(N434), .Z(n502) );
  CKBD1 U559 ( .I(N434), .Z(n501) );
  CKBD1 U560 ( .I(N434), .Z(n500) );
  CKBD1 U561 ( .I(N434), .Z(n499) );
  CKBD1 U562 ( .I(N434), .Z(n498) );
  CKBD1 U563 ( .I(N450), .Z(n382) );
  CKBD1 U564 ( .I(N450), .Z(n381) );
  CKBD1 U565 ( .I(N450), .Z(n380) );
  CKBD1 U566 ( .I(N450), .Z(n379) );
  CKBD1 U567 ( .I(N450), .Z(n378) );
  CKBD1 U568 ( .I(n582), .Z(n277) );
  CKBD1 U569 ( .I(n582), .Z(n276) );
  CKBD1 U570 ( .I(n582), .Z(n275) );
  CKBD1 U571 ( .I(n582), .Z(n274) );
  CKBD1 U572 ( .I(n582), .Z(n273) );
  CKBD1 U573 ( .I(N444), .Z(n427) );
  CKBD1 U574 ( .I(N444), .Z(n426) );
  CKBD1 U575 ( .I(N444), .Z(n425) );
  CKBD1 U576 ( .I(N444), .Z(n424) );
  CKBD1 U577 ( .I(N444), .Z(n423) );
  CKBD1 U578 ( .I(N460), .Z(n307) );
  CKBD1 U579 ( .I(N460), .Z(n306) );
  CKBD1 U580 ( .I(N460), .Z(n305) );
  CKBD1 U581 ( .I(N460), .Z(n304) );
  CKBD1 U582 ( .I(N460), .Z(n303) );
  CKBD1 U583 ( .I(n583), .Z(n292) );
  CKBD1 U584 ( .I(n583), .Z(n291) );
  CKBD1 U585 ( .I(n583), .Z(n290) );
  CKBD1 U586 ( .I(n583), .Z(n289) );
  CKBD1 U587 ( .I(n583), .Z(n288) );
  TIEH U588 ( .Z(RE) );
  TIEL U589 ( .ZN(WE) );
  NR2D0 U590 ( .A1(n533), .A2(n534), .ZN(n582) );
  NR2D0 U591 ( .A1(n534), .A2(n535), .ZN(n583) );
  CKND0 U592 ( .I(n536), .ZN(n585) );
  CKND2D0 U593 ( .A1(n584), .A2(op_done), .ZN(n537) );
  NR2D0 U594 ( .A1(n538), .A2(n545), .ZN(N460) );
  NR2D0 U595 ( .A1(n539), .A2(n545), .ZN(N458) );
  NR2D0 U596 ( .A1(n540), .A2(n545), .ZN(N456) );
  NR2D0 U597 ( .A1(n541), .A2(n545), .ZN(N454) );
  NR2D0 U598 ( .A1(n542), .A2(n545), .ZN(N452) );
  NR2D0 U599 ( .A1(n543), .A2(n545), .ZN(N450) );
  NR2D0 U600 ( .A1(n536), .A2(n545), .ZN(N448) );
  NR2D0 U601 ( .A1(n544), .A2(n545), .ZN(N446) );
  OR2D0 U602 ( .A1(n546), .A2(n534), .Z(n545) );
  NR2D0 U603 ( .A1(n538), .A2(n547), .ZN(N444) );
  NR2D0 U604 ( .A1(n539), .A2(n547), .ZN(N442) );
  NR2D0 U605 ( .A1(n540), .A2(n547), .ZN(N440) );
  NR2D0 U606 ( .A1(n541), .A2(n547), .ZN(N438) );
  NR2D0 U607 ( .A1(n542), .A2(n547), .ZN(N436) );
  NR2D0 U608 ( .A1(n543), .A2(n547), .ZN(N434) );
  NR2D0 U609 ( .A1(n536), .A2(n547), .ZN(N432) );
  NR2D0 U610 ( .A1(n544), .A2(n547), .ZN(N430) );
  OR2D0 U611 ( .A1(n548), .A2(n534), .Z(n547) );
  AOI21D0 U612 ( .A1(n549), .A2(n550), .B(n534), .ZN(N428) );
  CKND0 U613 ( .I(op_done), .ZN(n534) );
  INR2D0 U614 ( .A1(neuron_BAR[9]), .B1(n551), .ZN(N328) );
  XNR2D0 U615 ( .A1(neuron_BAR[9]), .A2(n551), .ZN(N327) );
  IND3D0 U616 ( .A1(n552), .B1(neuron_BAR[7]), .B2(neuron_BAR[8]), .ZN(n551)
         );
  XNR2D0 U617 ( .A1(n553), .A2(neuron_BAR[8]), .ZN(N326) );
  IND2D0 U618 ( .A1(n552), .B1(neuron_BAR[7]), .ZN(n553) );
  XNR2D0 U619 ( .A1(n552), .A2(neuron_BAR[7]), .ZN(N325) );
  AOI22D0 U620 ( .A1(n554), .A2(n555), .B1(n556), .B2(neuron_BAR[6]), .ZN(n552) );
  IND2D0 U621 ( .A1(n554), .B1(n549), .ZN(n556) );
  XOR3D0 U622 ( .A1(neuron_BAR[6]), .A2(n555), .A3(n554), .Z(N324) );
  MAOI222D0 U623 ( .A(n557), .B(n558), .C(n559), .ZN(n554) );
  CKND0 U624 ( .I(neuron_BAR[5]), .ZN(n557) );
  XOR3D0 U625 ( .A1(neuron_BAR[5]), .A2(n559), .A3(n558), .Z(N323) );
  AOI22D0 U626 ( .A1(n560), .A2(n561), .B1(n562), .B2(neuron_BAR[4]), .ZN(n558) );
  CKND2D0 U627 ( .A1(n563), .A2(n564), .ZN(n562) );
  CKND0 U628 ( .I(n563), .ZN(n561) );
  XOR3D0 U629 ( .A1(neuron_BAR[4]), .A2(n564), .A3(n563), .Z(N322) );
  IND3D0 U630 ( .A1(n565), .B1(neuron_BAR[2]), .B2(neuron_BAR[3]), .ZN(n563)
         );
  XNR2D0 U631 ( .A1(n566), .A2(neuron_BAR[3]), .ZN(N321) );
  IND2D0 U632 ( .A1(n565), .B1(neuron_BAR[2]), .ZN(n566) );
  XNR2D0 U633 ( .A1(n565), .A2(neuron_BAR[2]), .ZN(N320) );
  CKND0 U634 ( .I(n550), .ZN(N317) );
  NR2D0 U635 ( .A1(N315), .A2(\U3/U1/Z_5 ), .ZN(n550) );
  CKND0 U636 ( .I(n559), .ZN(\U3/U1/Z_5 ) );
  NR2D0 U637 ( .A1(n584), .A2(n567), .ZN(n559) );
  CKND0 U638 ( .I(n568), .ZN(n584) );
  IND2D0 U639 ( .A1(n567), .B1(n546), .ZN(N314) );
  IND2D0 U640 ( .A1(N315), .B1(n565), .ZN(N313) );
  NR2D0 U641 ( .A1(n567), .A2(n555), .ZN(n565) );
  CKND0 U642 ( .I(n549), .ZN(n555) );
  CKND2D0 U643 ( .A1(n533), .A2(n535), .ZN(n567) );
  CKND2D0 U644 ( .A1(n548), .A2(n546), .ZN(N315) );
  ND3D0 U645 ( .A1(n569), .A2(n570), .A3(n571), .ZN(n535) );
  ND3D0 U646 ( .A1(n572), .A2(mem_cur_state[0]), .A3(mem_cur_state[1]), .ZN(
        n568) );
  ND3D0 U647 ( .A1(n572), .A2(n569), .A3(mem_cur_state[1]), .ZN(n546) );
  CKND0 U648 ( .I(n560), .ZN(n564) );
  ND3D0 U649 ( .A1(n548), .A2(n533), .A3(n549), .ZN(n560) );
  ND3D0 U650 ( .A1(n571), .A2(n569), .A3(mem_cur_state[1]), .ZN(n549) );
  CKND0 U651 ( .I(mem_cur_state[0]), .ZN(n569) );
  ND3D0 U652 ( .A1(n571), .A2(n570), .A3(mem_cur_state[0]), .ZN(n533) );
  AN2D0 U653 ( .A1(mem_cur_state[3]), .A2(mem_cur_state[2]), .Z(n571) );
  ND3D0 U654 ( .A1(mem_cur_state[0]), .A2(n570), .A3(n572), .ZN(n548) );
  INR2D0 U655 ( .A1(mem_cur_state[3]), .B1(mem_cur_state[2]), .ZN(n572) );
  CKND0 U656 ( .I(mem_cur_state[1]), .ZN(n570) );
  NR4D0 U657 ( .A1(mem_cur_state[3]), .A2(mem_cur_state[2]), .A3(
        mem_cur_state[1]), .A4(mem_cur_state[0]), .ZN(N156) );
  ND3D0 U658 ( .A1(n542), .A2(n538), .A3(n573), .ZN(N124) );
  OAI211D0 U659 ( .A1(cur_state[0]), .A2(n574), .B(n541), .C(n573), .ZN(N123)
         );
  IND2D0 U660 ( .A1(N114), .B1(n574), .ZN(N122) );
  ND3D0 U661 ( .A1(n544), .A2(n540), .A3(n575), .ZN(N119) );
  ND3D0 U662 ( .A1(n540), .A2(n536), .A3(n573), .ZN(N118) );
  CKND2D0 U663 ( .A1(n575), .A2(n576), .ZN(N117) );
  ND3D0 U664 ( .A1(n540), .A2(n576), .A3(n541), .ZN(N116) );
  ND3D0 U665 ( .A1(n544), .A2(n541), .A3(n573), .ZN(N115) );
  AN2D0 U666 ( .A1(n539), .A2(n543), .Z(n573) );
  IND4D0 U667 ( .A1(N125), .B1(n538), .B2(n539), .B3(n576), .ZN(N114) );
  CKND0 U668 ( .I(N121), .ZN(n576) );
  CKND2D0 U669 ( .A1(n536), .A2(n544), .ZN(N121) );
  ND4D0 U670 ( .A1(cur_state[3]), .A2(n577), .A3(n578), .A4(n579), .ZN(n544)
         );
  ND3D0 U671 ( .A1(cur_state[0]), .A2(n580), .A3(cur_state[1]), .ZN(n536) );
  ND4D0 U672 ( .A1(cur_state[1]), .A2(n577), .A3(n579), .A4(n581), .ZN(n539)
         );
  IND2D0 U673 ( .A1(n574), .B1(cur_state[0]), .ZN(n538) );
  ND3D0 U674 ( .A1(n579), .A2(n581), .A3(n578), .ZN(n574) );
  IND2D0 U675 ( .A1(N120), .B1(n540), .ZN(N125) );
  ND4D0 U676 ( .A1(cur_state[1]), .A2(cur_state[0]), .A3(n579), .A4(n581), 
        .ZN(n540) );
  CKND0 U677 ( .I(cur_state[3]), .ZN(n581) );
  CKND2D0 U678 ( .A1(n575), .A2(n541), .ZN(N120) );
  ND3D0 U679 ( .A1(n577), .A2(n578), .A3(n580), .ZN(n541) );
  AN2D0 U680 ( .A1(n542), .A2(n543), .Z(n575) );
  ND3D0 U681 ( .A1(n580), .A2(n577), .A3(cur_state[1]), .ZN(n543) );
  CKND0 U682 ( .I(cur_state[0]), .ZN(n577) );
  ND3D0 U683 ( .A1(n580), .A2(n578), .A3(cur_state[0]), .ZN(n542) );
  CKND0 U684 ( .I(cur_state[1]), .ZN(n578) );
  NR2D0 U685 ( .A1(n579), .A2(cur_state[3]), .ZN(n580) );
  CKND0 U686 ( .I(cur_state[2]), .ZN(n579) );
endmodule

