
module fma_lza ( mantissa_ab, mantissa_c, exp_ab_greater, exp_ab_less, sign_ab, 
        sign_c, fma_byp, adder_start, mantissa_shift, lza_done );
  input [21:0] mantissa_ab;
  input [21:0] mantissa_c;
  output [4:0] mantissa_shift;
  input exp_ab_greater, exp_ab_less, sign_ab, sign_c, fma_byp, adder_start;
  output lza_done;
  wire   adder_start, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167;
  assign lza_done = adder_start;

  NR3D2 U3 ( .A1(n63), .A2(n1), .A3(n64), .ZN(mantissa_shift[1]) );
  XNR2D1 U4 ( .A1(n62), .A2(n61), .ZN(n63) );
  NR2D3 U5 ( .A1(n1), .A2(n2), .ZN(mantissa_shift[4]) );
  NR2D3 U6 ( .A1(n1), .A2(n15), .ZN(mantissa_shift[3]) );
  NR2D3 U7 ( .A1(n94), .A2(n1), .ZN(mantissa_shift[0]) );
  NR2D3 U8 ( .A1(n1), .A2(n31), .ZN(mantissa_shift[2]) );
  CKXOR2D0 U9 ( .A1(n3), .A2(n4), .Z(n2) );
  MUX2ND0 U10 ( .I0(n5), .I1(n6), .S(n7), .ZN(n4) );
  CKND2D0 U11 ( .A1(n8), .A2(n9), .ZN(n6) );
  CKND2D0 U12 ( .A1(n10), .A2(n11), .ZN(n5) );
  AOI21D0 U13 ( .A1(n12), .A2(n13), .B(n14), .ZN(n3) );
  XNR3D0 U14 ( .A1(n12), .A2(n14), .A3(n13), .ZN(n15) );
  MUX2D0 U15 ( .I0(n16), .I1(n17), .S(sign_c), .Z(n13) );
  XNR2D0 U16 ( .A1(n11), .A2(n10), .ZN(n17) );
  AOI21D0 U17 ( .A1(n18), .A2(n10), .B(n19), .ZN(n11) );
  XNR2D0 U18 ( .A1(n9), .A2(n8), .ZN(n16) );
  AOI21D0 U19 ( .A1(n20), .A2(n8), .B(n21), .ZN(n9) );
  OAI21D0 U20 ( .A1(n22), .A2(n23), .B(n24), .ZN(n14) );
  MUX2D0 U21 ( .I0(n25), .I1(n26), .S(sign_c), .Z(n12) );
  CKND2D0 U22 ( .A1(n27), .A2(n28), .ZN(n26) );
  CKND2D0 U23 ( .A1(n29), .A2(n30), .ZN(n25) );
  CKXOR2D0 U24 ( .A1(n32), .A2(n23), .Z(n31) );
  MUX2ND0 U25 ( .I0(n33), .I1(n34), .S(n7), .ZN(n23) );
  XNR2D0 U26 ( .A1(n30), .A2(n35), .ZN(n34) );
  OA21D0 U27 ( .A1(n36), .A2(n37), .B(n29), .Z(n35) );
  NR2D0 U28 ( .A1(n38), .A2(n39), .ZN(n29) );
  XNR2D0 U29 ( .A1(n28), .A2(n40), .ZN(n33) );
  OA21D0 U30 ( .A1(n41), .A2(n42), .B(n27), .Z(n40) );
  NR2D0 U31 ( .A1(n43), .A2(n44), .ZN(n27) );
  INR2D0 U32 ( .A1(n24), .B1(n22), .ZN(n32) );
  MUX2ND0 U33 ( .I0(n45), .I1(n46), .S(n7), .ZN(n22) );
  XOR3D0 U34 ( .A1(n8), .A2(n20), .A3(n21), .Z(n46) );
  AO21D0 U35 ( .A1(n47), .A2(n48), .B(n49), .Z(n21) );
  CKND2D0 U36 ( .A1(n50), .A2(n51), .ZN(n20) );
  NR2D0 U37 ( .A1(n52), .A2(n53), .ZN(n8) );
  XOR3D0 U38 ( .A1(n10), .A2(n18), .A3(n19), .Z(n45) );
  AO21D0 U39 ( .A1(n54), .A2(n55), .B(n56), .Z(n19) );
  CKND2D0 U40 ( .A1(n57), .A2(n58), .ZN(n18) );
  NR2D0 U41 ( .A1(n59), .A2(n60), .ZN(n10) );
  INR2D0 U42 ( .A1(n61), .B1(n62), .ZN(n24) );
  MUX2ND0 U43 ( .I0(n65), .I1(n66), .S(n7), .ZN(n64) );
  CKND2D0 U44 ( .A1(n47), .A2(n67), .ZN(n66) );
  CKXOR2D0 U45 ( .A1(n49), .A2(n48), .Z(n67) );
  AN2D0 U46 ( .A1(n68), .A2(n69), .Z(n48) );
  XNR2D0 U47 ( .A1(n51), .A2(n50), .ZN(n68) );
  INR2D0 U48 ( .A1(n70), .B1(n71), .ZN(n49) );
  CKXOR2D0 U49 ( .A1(n72), .A2(n53), .Z(n47) );
  NR2D0 U50 ( .A1(n73), .A2(n52), .ZN(n72) );
  NR2D0 U51 ( .A1(n74), .A2(n75), .ZN(n52) );
  CKND2D0 U52 ( .A1(n54), .A2(n76), .ZN(n65) );
  CKXOR2D0 U53 ( .A1(n55), .A2(n56), .Z(n76) );
  AN2D0 U54 ( .A1(n77), .A2(n78), .Z(n55) );
  XNR2D0 U55 ( .A1(n58), .A2(n57), .ZN(n77) );
  XNR2D0 U56 ( .A1(n59), .A2(n60), .ZN(n54) );
  MUX2ND0 U57 ( .I0(n79), .I1(n80), .S(n7), .ZN(n61) );
  INR3D0 U58 ( .A1(n30), .B1(n81), .B2(n82), .ZN(n80) );
  XNR2D0 U59 ( .A1(n36), .A2(n83), .ZN(n81) );
  CKND2D0 U60 ( .A1(n84), .A2(n85), .ZN(n30) );
  XNR2D0 U61 ( .A1(n86), .A2(n87), .ZN(n84) );
  INR3D0 U62 ( .A1(n28), .B1(n88), .B2(n89), .ZN(n79) );
  CKXOR2D0 U63 ( .A1(n41), .A2(n42), .Z(n88) );
  CKND2D0 U64 ( .A1(n90), .A2(n91), .ZN(n28) );
  XNR2D0 U65 ( .A1(n44), .A2(n43), .ZN(n90) );
  INR2D0 U66 ( .A1(n92), .B1(n93), .ZN(n62) );
  OR2D0 U67 ( .A1(fma_byp), .A2(sign_ab), .Z(n1) );
  CKXOR2D0 U68 ( .A1(n93), .A2(n92), .Z(n94) );
  OAI31D0 U69 ( .A1(n7), .A2(n95), .A3(n56), .B(n96), .ZN(n92) );
  CKXOR2D0 U70 ( .A1(n70), .A2(n71), .Z(n96) );
  CKND2D0 U71 ( .A1(n97), .A2(n50), .ZN(n71) );
  XNR2D0 U72 ( .A1(n98), .A2(n99), .ZN(n50) );
  NR2D0 U73 ( .A1(n100), .A2(n101), .ZN(n98) );
  OAI21D0 U74 ( .A1(n69), .A2(n102), .B(n103), .ZN(n97) );
  CKXOR2D0 U75 ( .A1(n74), .A2(n75), .Z(n70) );
  ND4D0 U76 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(n75) );
  NR4D0 U77 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(n107) );
  AO33D0 U78 ( .A1(n112), .A2(mantissa_ab[20]), .A3(mantissa_c[20]), .B1(
        mantissa_c[19]), .B2(n113), .B3(mantissa_ab[19]), .Z(n111) );
  AO31D0 U79 ( .A1(n114), .A2(mantissa_ab[18]), .A3(mantissa_c[18]), .B(n115), 
        .Z(n110) );
  AO33D0 U80 ( .A1(mantissa_ab[16]), .A2(n37), .A3(mantissa_c[16]), .B1(
        mantissa_c[17]), .B2(mantissa_ab[17]), .B3(n116), .Z(n115) );
  OAI31D0 U81 ( .A1(n117), .A2(n118), .A3(n119), .B(n120), .ZN(n109) );
  AOI33D0 U82 ( .A1(mantissa_ab[13]), .A2(n85), .A3(mantissa_c[13]), .B1(
        mantissa_c[14]), .B2(mantissa_ab[14]), .B3(n121), .ZN(n120) );
  AO31D0 U83 ( .A1(n122), .A2(mantissa_ab[12]), .A3(mantissa_c[12]), .B(n123), 
        .Z(n108) );
  AO33D0 U84 ( .A1(mantissa_ab[10]), .A2(n39), .A3(mantissa_c[10]), .B1(
        mantissa_c[11]), .B2(mantissa_ab[11]), .B3(n124), .Z(n123) );
  NR4D0 U85 ( .A1(n125), .A2(n126), .A3(n127), .A4(n73), .ZN(n106) );
  INR3D0 U86 ( .A1(n128), .B1(mantissa_ab[0]), .B2(mantissa_c[0]), .ZN(n73) );
  AN3D0 U87 ( .A1(n128), .A2(mantissa_ab[0]), .A3(mantissa_c[0]), .Z(n126) );
  AO31D0 U88 ( .A1(n100), .A2(mantissa_ab[3]), .A3(mantissa_c[3]), .B(n129), 
        .Z(n125) );
  AO33D0 U89 ( .A1(mantissa_ab[1]), .A2(n53), .A3(mantissa_c[1]), .B1(
        mantissa_c[2]), .B2(mantissa_ab[2]), .B3(n130), .Z(n129) );
  AOI31D0 U90 ( .A1(mantissa_c[6]), .A2(mantissa_ab[6]), .A3(n131), .B(n132), 
        .ZN(n105) );
  AO33D0 U91 ( .A1(n133), .A2(mantissa_ab[5]), .A3(mantissa_c[5]), .B1(
        mantissa_c[4]), .B2(n99), .B3(mantissa_ab[4]), .Z(n132) );
  AOI31D0 U92 ( .A1(mantissa_ab[9]), .A2(n134), .A3(mantissa_c[9]), .B(n135), 
        .ZN(n104) );
  AO33D0 U93 ( .A1(n136), .A2(mantissa_ab[8]), .A3(mantissa_c[8]), .B1(
        mantissa_c[7]), .B2(n69), .B3(mantissa_ab[7]), .Z(n135) );
  AOI21D0 U94 ( .A1(n137), .A2(n130), .B(n128), .ZN(n74) );
  NR3D0 U95 ( .A1(mantissa_ab[1]), .A2(mantissa_c[1]), .A3(n137), .ZN(n128) );
  CKND0 U96 ( .I(n53), .ZN(n137) );
  INR3D0 U97 ( .A1(n130), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n53) );
  INR3D0 U98 ( .A1(n100), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n130)
         );
  NR3D0 U99 ( .A1(mantissa_ab[4]), .A2(mantissa_c[4]), .A3(n51), .ZN(n100) );
  CKND0 U100 ( .I(n99), .ZN(n51) );
  NR3D0 U101 ( .A1(mantissa_ab[5]), .A2(mantissa_c[5]), .A3(n101), .ZN(n99) );
  CKND0 U102 ( .I(n133), .ZN(n101) );
  NR3D0 U103 ( .A1(mantissa_ab[6]), .A2(mantissa_c[6]), .A3(n103), .ZN(n133)
         );
  CKND0 U104 ( .I(n131), .ZN(n103) );
  INR3D0 U105 ( .A1(n69), .B1(mantissa_ab[7]), .B2(mantissa_c[7]), .ZN(n131)
         );
  NR3D0 U106 ( .A1(mantissa_ab[8]), .A2(mantissa_c[8]), .A3(n102), .ZN(n69) );
  CKND0 U107 ( .I(n136), .ZN(n102) );
  INR3D0 U108 ( .A1(n134), .B1(mantissa_ab[9]), .B2(mantissa_c[9]), .ZN(n136)
         );
  OA21D0 U109 ( .A1(n138), .A2(n139), .B(n57), .Z(n56) );
  OA21D0 U110 ( .A1(n140), .A2(n141), .B(n142), .Z(n57) );
  NR2D0 U111 ( .A1(n78), .A2(n143), .ZN(n139) );
  AOI31D0 U112 ( .A1(mantissa_ab[0]), .A2(n144), .A3(mantissa_c[0]), .B(n145), 
        .ZN(n95) );
  CKND0 U113 ( .I(n60), .ZN(n145) );
  OAI21D0 U114 ( .A1(n59), .A2(n146), .B(n147), .ZN(n60) );
  CKND0 U115 ( .I(n147), .ZN(n144) );
  ND3D0 U116 ( .A1(mantissa_ab[1]), .A2(n59), .A3(mantissa_c[1]), .ZN(n147) );
  CKND0 U117 ( .I(n148), .ZN(n59) );
  IND3D0 U118 ( .A1(n146), .B1(mantissa_ab[2]), .B2(mantissa_c[2]), .ZN(n148)
         );
  IND3D0 U119 ( .A1(n142), .B1(mantissa_ab[3]), .B2(mantissa_c[3]), .ZN(n146)
         );
  ND3D0 U120 ( .A1(mantissa_ab[4]), .A2(n140), .A3(mantissa_c[4]), .ZN(n142)
         );
  CKND0 U121 ( .I(n58), .ZN(n140) );
  IND3D0 U122 ( .A1(n141), .B1(mantissa_ab[5]), .B2(mantissa_c[5]), .ZN(n58)
         );
  ND3D0 U123 ( .A1(mantissa_ab[6]), .A2(n138), .A3(mantissa_c[6]), .ZN(n141)
         );
  AN3D0 U124 ( .A1(mantissa_ab[7]), .A2(n78), .A3(mantissa_c[7]), .Z(n138) );
  AN3D0 U125 ( .A1(n149), .A2(mantissa_ab[8]), .A3(mantissa_c[8]), .Z(n78) );
  CKND0 U126 ( .I(n143), .ZN(n149) );
  IND3D0 U127 ( .A1(n150), .B1(mantissa_ab[9]), .B2(mantissa_c[9]), .ZN(n143)
         );
  MUX2ND0 U128 ( .I0(n151), .I1(n152), .S(n7), .ZN(n93) );
  CKND0 U129 ( .I(sign_c), .ZN(n7) );
  OAI22D0 U130 ( .A1(n36), .A2(n153), .B1(n38), .B2(n154), .ZN(n152) );
  AOI21D0 U131 ( .A1(n121), .A2(n155), .B(n122), .ZN(n154) );
  CKND0 U132 ( .I(n87), .ZN(n38) );
  AOI21D0 U133 ( .A1(n86), .A2(n124), .B(n134), .ZN(n87) );
  NR3D0 U134 ( .A1(mantissa_ab[10]), .A2(mantissa_c[10]), .A3(n86), .ZN(n134)
         );
  CKND0 U135 ( .I(n39), .ZN(n86) );
  INR3D0 U136 ( .A1(n124), .B1(mantissa_ab[11]), .B2(mantissa_c[11]), .ZN(n39)
         );
  INR3D0 U137 ( .A1(n122), .B1(mantissa_ab[12]), .B2(mantissa_c[12]), .ZN(n124) );
  NR3D0 U138 ( .A1(mantissa_ab[13]), .A2(mantissa_c[13]), .A3(n155), .ZN(n122)
         );
  CKND0 U139 ( .I(n85), .ZN(n155) );
  INR3D0 U140 ( .A1(n121), .B1(mantissa_ab[14]), .B2(mantissa_c[14]), .ZN(n85)
         );
  NR3D0 U141 ( .A1(mantissa_ab[15]), .A2(mantissa_c[15]), .A3(n117), .ZN(n121)
         );
  AOI21D0 U142 ( .A1(n112), .A2(n82), .B(n114), .ZN(n153) );
  IOA21D0 U143 ( .A1(n83), .A2(n116), .B(n117), .ZN(n36) );
  OR3D0 U144 ( .A1(mantissa_ab[16]), .A2(mantissa_c[16]), .A3(n83), .Z(n117)
         );
  CKND0 U145 ( .I(n37), .ZN(n83) );
  INR3D0 U146 ( .A1(n116), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n37)
         );
  INR3D0 U147 ( .A1(n114), .B1(mantissa_ab[18]), .B2(mantissa_c[18]), .ZN(n116) );
  NR3D0 U148 ( .A1(mantissa_ab[19]), .A2(mantissa_c[19]), .A3(n82), .ZN(n114)
         );
  CKND0 U149 ( .I(n113), .ZN(n82) );
  INR3D0 U150 ( .A1(n112), .B1(mantissa_ab[20]), .B2(mantissa_c[20]), .ZN(n113) );
  NR2D0 U151 ( .A1(mantissa_ab[21]), .A2(mantissa_c[21]), .ZN(n112) );
  OAI22D0 U152 ( .A1(n41), .A2(n156), .B1(n43), .B2(n157), .ZN(n151) );
  AOI21D0 U153 ( .A1(n158), .A2(n159), .B(n160), .ZN(n157) );
  OAI21D0 U154 ( .A1(n44), .A2(n161), .B(n150), .ZN(n43) );
  ND3D0 U155 ( .A1(mantissa_ab[10]), .A2(n44), .A3(mantissa_c[10]), .ZN(n150)
         );
  AN3D0 U156 ( .A1(n162), .A2(mantissa_ab[11]), .A3(mantissa_c[11]), .Z(n44)
         );
  CKND0 U157 ( .I(n161), .ZN(n162) );
  ND3D0 U158 ( .A1(mantissa_ab[12]), .A2(n160), .A3(mantissa_c[12]), .ZN(n161)
         );
  AN3D0 U159 ( .A1(mantissa_ab[13]), .A2(n91), .A3(mantissa_c[13]), .Z(n160)
         );
  CKND0 U160 ( .I(n159), .ZN(n91) );
  ND3D0 U161 ( .A1(mantissa_ab[14]), .A2(n158), .A3(mantissa_c[14]), .ZN(n159)
         );
  NR3D0 U162 ( .A1(n118), .A2(n163), .A3(n119), .ZN(n158) );
  CKND0 U163 ( .I(mantissa_c[15]), .ZN(n119) );
  CKND0 U164 ( .I(mantissa_ab[15]), .ZN(n118) );
  AOI21D0 U165 ( .A1(n127), .A2(n89), .B(n164), .ZN(n156) );
  OAI21D0 U166 ( .A1(n42), .A2(n165), .B(n163), .ZN(n41) );
  ND3D0 U167 ( .A1(mantissa_ab[16]), .A2(n42), .A3(mantissa_c[16]), .ZN(n163)
         );
  CKND0 U168 ( .I(n166), .ZN(n42) );
  IND3D0 U169 ( .A1(n165), .B1(mantissa_ab[17]), .B2(mantissa_c[17]), .ZN(n166) );
  ND3D0 U170 ( .A1(mantissa_ab[18]), .A2(n164), .A3(mantissa_c[18]), .ZN(n165)
         );
  CKND0 U171 ( .I(n167), .ZN(n164) );
  IND3D0 U172 ( .A1(n89), .B1(mantissa_ab[19]), .B2(mantissa_c[19]), .ZN(n167)
         );
  ND3D0 U173 ( .A1(mantissa_ab[20]), .A2(n127), .A3(mantissa_c[20]), .ZN(n89)
         );
  AN2D0 U174 ( .A1(mantissa_c[21]), .A2(mantissa_ab[21]), .Z(n127) );
endmodule


module fma_aligner_adder_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [20:0] A;
  input [4:0] SH;
  output [20:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  INVD1 U3 ( .I(n61), .ZN(n14) );
  INVD1 U4 ( .I(n53), .ZN(n22) );
  INVD1 U5 ( .I(n52), .ZN(n23) );
  INVD1 U6 ( .I(n47), .ZN(n15) );
  INVD1 U7 ( .I(n81), .ZN(n20) );
  INVD1 U8 ( .I(n58), .ZN(n3) );
  INVD1 U9 ( .I(n80), .ZN(n21) );
  INVD1 U10 ( .I(n27), .ZN(n1) );
  INVD1 U11 ( .I(n37), .ZN(n17) );
  INVD1 U12 ( .I(n25), .ZN(n8) );
  INVD1 U13 ( .I(n59), .ZN(n7) );
  INVD1 U14 ( .I(n51), .ZN(n6) );
  INVD1 U15 ( .I(n70), .ZN(n5) );
  INVD1 U16 ( .I(n50), .ZN(n2) );
  INVD1 U17 ( .I(n36), .ZN(n16) );
  INVD1 U18 ( .I(n29), .ZN(n9) );
  INVD1 U19 ( .I(n30), .ZN(n4) );
  INVD1 U20 ( .I(SH[2]), .ZN(n19) );
  INVD1 U21 ( .I(A[3]), .ZN(n11) );
  INVD1 U22 ( .I(A[2]), .ZN(n12) );
  INVD1 U23 ( .I(SH[3]), .ZN(n18) );
  INVD1 U24 ( .I(SH[0]), .ZN(n24) );
  INVD1 U25 ( .I(A[4]), .ZN(n10) );
  INVD1 U26 ( .I(A[1]), .ZN(n13) );
  OAI222D0 U27 ( .A1(n25), .A2(n26), .B1(n27), .B2(n17), .C1(n28), .C2(n15), 
        .ZN(B[9]) );
  OAI222D0 U28 ( .A1(n29), .A2(n26), .B1(n30), .B2(n31), .C1(n32), .C2(n15), 
        .ZN(B[8]) );
  OAI221D0 U29 ( .A1(n33), .A2(n26), .B1(n34), .B2(n15), .C(n35), .ZN(B[7]) );
  AOI22D0 U30 ( .A1(n36), .A2(n2), .B1(n37), .B2(n6), .ZN(n35) );
  OAI221D0 U31 ( .A1(n38), .A2(n26), .B1(n39), .B2(n15), .C(n40), .ZN(B[6]) );
  AOI22D0 U32 ( .A1(n36), .A2(n3), .B1(n37), .B2(n7), .ZN(n40) );
  OAI221D0 U33 ( .A1(n28), .A2(n26), .B1(n41), .B2(n15), .C(n42), .ZN(B[5]) );
  AOI22D0 U34 ( .A1(n36), .A2(n1), .B1(n37), .B2(n8), .ZN(n42) );
  OAI221D0 U35 ( .A1(n32), .A2(n26), .B1(n43), .B2(n15), .C(n44), .ZN(B[4]) );
  AOI222D0 U36 ( .A1(n37), .A2(n9), .B1(n45), .B2(n14), .C1(n36), .C2(n5), 
        .ZN(n44) );
  OAI221D0 U37 ( .A1(n33), .A2(n17), .B1(n34), .B2(n26), .C(n46), .ZN(B[3]) );
  AOI222D0 U38 ( .A1(n36), .A2(n6), .B1(n45), .B2(n2), .C1(n47), .C2(n48), 
        .ZN(n46) );
  OAI221D0 U39 ( .A1(n23), .A2(n10), .B1(n22), .B2(n11), .C(n49), .ZN(n48) );
  AOI22D0 U40 ( .A1(A[6]), .A2(n21), .B1(A[5]), .B2(n20), .ZN(n49) );
  AOI221D0 U41 ( .A1(n52), .A2(A[8]), .B1(n53), .B2(A[7]), .C(n54), .ZN(n34)
         );
  AO22D0 U42 ( .A1(A[10]), .A2(n21), .B1(A[9]), .B2(n20), .Z(n54) );
  OAI221D0 U43 ( .A1(n38), .A2(n17), .B1(n39), .B2(n26), .C(n55), .ZN(B[2]) );
  AOI222D0 U44 ( .A1(n36), .A2(n7), .B1(n45), .B2(n3), .C1(n47), .C2(n56), 
        .ZN(n55) );
  OAI221D0 U45 ( .A1(n23), .A2(n11), .B1(n22), .B2(n12), .C(n57), .ZN(n56) );
  AOI22D0 U46 ( .A1(A[5]), .A2(n21), .B1(A[4]), .B2(n20), .ZN(n57) );
  AOI221D0 U47 ( .A1(n52), .A2(A[7]), .B1(n53), .B2(A[6]), .C(n60), .ZN(n39)
         );
  AO22D0 U48 ( .A1(A[9]), .A2(n21), .B1(A[8]), .B2(n20), .Z(n60) );
  NR2D0 U49 ( .A1(n15), .A2(n61), .ZN(B[20]) );
  OAI221D0 U50 ( .A1(n28), .A2(n17), .B1(n41), .B2(n26), .C(n62), .ZN(B[1]) );
  AOI222D0 U51 ( .A1(n36), .A2(n8), .B1(n45), .B2(n1), .C1(n47), .C2(n63), 
        .ZN(n62) );
  OAI221D0 U52 ( .A1(n23), .A2(n12), .B1(n22), .B2(n13), .C(n64), .ZN(n63) );
  AOI22D0 U53 ( .A1(A[4]), .A2(n21), .B1(A[3]), .B2(n20), .ZN(n64) );
  AN3D0 U54 ( .A1(SH[4]), .A2(n19), .A3(n18), .Z(n45) );
  AOI221D0 U55 ( .A1(n52), .A2(A[6]), .B1(n53), .B2(A[5]), .C(n65), .ZN(n41)
         );
  AO22D0 U56 ( .A1(A[8]), .A2(n21), .B1(A[7]), .B2(n20), .Z(n65) );
  AOI221D0 U57 ( .A1(n52), .A2(A[10]), .B1(n53), .B2(A[9]), .C(n66), .ZN(n28)
         );
  AO22D0 U58 ( .A1(A[12]), .A2(n21), .B1(A[11]), .B2(n20), .Z(n66) );
  NR2D0 U59 ( .A1(n50), .A2(n15), .ZN(B[19]) );
  NR2D0 U60 ( .A1(n58), .A2(n15), .ZN(B[18]) );
  NR2D0 U61 ( .A1(n27), .A2(n15), .ZN(B[17]) );
  NR2D0 U62 ( .A1(n30), .A2(n67), .ZN(B[16]) );
  OAI22D0 U63 ( .A1(n51), .A2(n15), .B1(n50), .B2(n26), .ZN(B[15]) );
  OAI22D0 U64 ( .A1(n59), .A2(n15), .B1(n58), .B2(n26), .ZN(B[14]) );
  OAI22D0 U65 ( .A1(n25), .A2(n15), .B1(n27), .B2(n26), .ZN(B[13]) );
  AOI221D0 U66 ( .A1(n52), .A2(A[18]), .B1(n53), .B2(A[17]), .C(n68), .ZN(n27)
         );
  AO22D0 U67 ( .A1(A[20]), .A2(n21), .B1(A[19]), .B2(n20), .Z(n68) );
  AOI221D0 U68 ( .A1(n52), .A2(A[14]), .B1(n53), .B2(A[13]), .C(n69), .ZN(n25)
         );
  AO22D0 U69 ( .A1(A[16]), .A2(n21), .B1(A[15]), .B2(n20), .Z(n69) );
  OAI222D0 U70 ( .A1(n70), .A2(n26), .B1(n17), .B2(n61), .C1(n29), .C2(n15), 
        .ZN(B[12]) );
  OAI222D0 U71 ( .A1(n51), .A2(n26), .B1(n50), .B2(n17), .C1(n33), .C2(n15), 
        .ZN(B[11]) );
  AOI221D0 U72 ( .A1(n52), .A2(A[12]), .B1(n53), .B2(A[11]), .C(n71), .ZN(n33)
         );
  AO22D0 U73 ( .A1(A[14]), .A2(n21), .B1(A[13]), .B2(n20), .Z(n71) );
  AOI22D0 U74 ( .A1(A[19]), .A2(n53), .B1(A[20]), .B2(n52), .ZN(n50) );
  AOI221D0 U75 ( .A1(n52), .A2(A[16]), .B1(n53), .B2(A[15]), .C(n72), .ZN(n51)
         );
  AO22D0 U76 ( .A1(A[18]), .A2(n21), .B1(A[17]), .B2(n20), .Z(n72) );
  OAI222D0 U77 ( .A1(n59), .A2(n26), .B1(n58), .B2(n17), .C1(n38), .C2(n15), 
        .ZN(B[10]) );
  AOI221D0 U78 ( .A1(n52), .A2(A[11]), .B1(n53), .B2(A[10]), .C(n73), .ZN(n38)
         );
  AO22D0 U79 ( .A1(A[13]), .A2(n21), .B1(A[12]), .B2(n20), .Z(n73) );
  AOI222D0 U80 ( .A1(A[19]), .A2(n52), .B1(A[20]), .B2(n20), .C1(A[18]), .C2(
        n53), .ZN(n58) );
  AOI221D0 U81 ( .A1(n52), .A2(A[15]), .B1(n53), .B2(A[14]), .C(n74), .ZN(n59)
         );
  AO22D0 U82 ( .A1(A[17]), .A2(n21), .B1(A[16]), .B2(n20), .Z(n74) );
  OAI211D0 U83 ( .A1(n29), .A2(n16), .B(n75), .C(n76), .ZN(B[0]) );
  OA22D0 U84 ( .A1(n17), .A2(n32), .B1(n26), .B2(n43), .Z(n76) );
  AOI221D0 U85 ( .A1(n52), .A2(A[5]), .B1(n53), .B2(A[4]), .C(n77), .ZN(n43)
         );
  AO22D0 U86 ( .A1(A[7]), .A2(n21), .B1(A[6]), .B2(n20), .Z(n77) );
  IND2D0 U87 ( .A1(n67), .B1(SH[2]), .ZN(n26) );
  AOI221D0 U88 ( .A1(n52), .A2(A[9]), .B1(n53), .B2(A[8]), .C(n78), .ZN(n32)
         );
  AO22D0 U89 ( .A1(A[11]), .A2(n21), .B1(A[10]), .B2(n20), .Z(n78) );
  NR2D0 U90 ( .A1(n31), .A2(SH[2]), .ZN(n37) );
  AOI32D0 U91 ( .A1(n4), .A2(n18), .A3(SH[4]), .B1(n47), .B2(n79), .ZN(n75) );
  OAI221D0 U92 ( .A1(n80), .A2(n11), .B1(n81), .B2(n12), .C(n82), .ZN(n79) );
  AOI22D0 U93 ( .A1(A[1]), .A2(n52), .B1(A[0]), .B2(n53), .ZN(n82) );
  NR2D0 U94 ( .A1(n67), .A2(SH[2]), .ZN(n47) );
  OR2D0 U95 ( .A1(SH[4]), .A2(SH[3]), .Z(n67) );
  MUX2ND0 U96 ( .I0(n14), .I1(n5), .S(n19), .ZN(n30) );
  AOI221D0 U97 ( .A1(n52), .A2(A[17]), .B1(n53), .B2(A[16]), .C(n83), .ZN(n70)
         );
  AO22D0 U98 ( .A1(A[19]), .A2(n21), .B1(A[18]), .B2(n20), .Z(n83) );
  CKND2D0 U99 ( .A1(n53), .A2(A[20]), .ZN(n61) );
  NR2D0 U100 ( .A1(n19), .A2(n31), .ZN(n36) );
  OR2D0 U101 ( .A1(SH[4]), .A2(n18), .Z(n31) );
  AOI221D0 U102 ( .A1(n52), .A2(A[13]), .B1(n53), .B2(A[12]), .C(n84), .ZN(n29) );
  AO22D0 U103 ( .A1(A[15]), .A2(n21), .B1(A[14]), .B2(n20), .Z(n84) );
  CKND2D0 U104 ( .A1(SH[1]), .A2(n24), .ZN(n81) );
  CKND2D0 U105 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  NR2D0 U106 ( .A1(SH[0]), .A2(SH[1]), .ZN(n53) );
  NR2D0 U107 ( .A1(n24), .A2(SH[1]), .ZN(n52) );
endmodule


module fma_aligner_adder ( mantissa_ab, exp_ab, sign_ab, c, exp_diff, 
        exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start, 
        mantissa_ab_c, exp_ab_c, sign_ab_c, mantissa_shift, adder_done );
  input [19:0] mantissa_ab;
  input [4:0] exp_ab;
  input [15:0] c;
  input [4:0] exp_diff;
  output [21:0] mantissa_ab_c;
  output [4:0] exp_ab_c;
  output [4:0] mantissa_shift;
  input sign_ab, exp_ab_greater, exp_ab_less, fma_byp, add_byp, adder_start;
  output sign_ab_c, adder_done;
  wire   n1147, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N800, n11, n535, n536,
         n537, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145;
  wire   [21:0] comp_mantissa_ab;
  wire   [21:0] comp_mantissa_c;

  fma_lza fma_lza_i ( .mantissa_ab(comp_mantissa_ab), .mantissa_c(
        comp_mantissa_c), .exp_ab_greater(exp_ab_greater), .exp_ab_less(
        exp_ab_less), .sign_ab(sign_ab), .sign_c(c[15]), .fma_byp(fma_byp), 
        .adder_start(adder_start), .mantissa_shift(mantissa_shift), .lza_done(
        adder_done) );
  fma_aligner_adder_DW_rash_0 srl_62 ( .A({N800, mantissa_ab}), .DATA_TC(n11), 
        .SH(exp_diff), .SH_TC(n11), .B({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45}) );
  OA21D1 U600 ( .A1(n563), .A2(n593), .B(n703), .Z(n535) );
  OA21D1 U601 ( .A1(n558), .A2(n593), .B(n671), .Z(n536) );
  OA21D1 U602 ( .A1(n627), .A2(n593), .B(n628), .Z(n537) );
  MUX2ND2 U603 ( .I0(n588), .I1(n589), .S(n590), .ZN(mantissa_ab_c[8]) );
  INVD2 U604 ( .I(n537), .ZN(mantissa_ab_c[20]) );
  INVD2 U605 ( .I(n536), .ZN(mantissa_ab_c[18]) );
  INVD2 U606 ( .I(n535), .ZN(mantissa_ab_c[16]) );
  OAI21D4 U607 ( .A1(n564), .A2(n593), .B(n714), .ZN(mantissa_ab_c[15]) );
  MUX2ND2 U608 ( .I0(n595), .I1(n596), .S(n597), .ZN(mantissa_ab_c[7]) );
  IAO21D1 U609 ( .A1(n598), .A2(fma_byp), .B(n594), .ZN(n595) );
  OAI21D4 U610 ( .A1(n572), .A2(n593), .B(n743), .ZN(mantissa_ab_c[13]) );
  MUX2ND2 U611 ( .I0(n613), .I1(n614), .S(n615), .ZN(mantissa_ab_c[3]) );
  ND2D1 U612 ( .A1(n583), .A2(n616), .ZN(n613) );
  OAI21D4 U613 ( .A1(n652), .A2(n593), .B(n653), .ZN(mantissa_ab_c[19]) );
  MUX2ND2 U614 ( .I0(n599), .I1(n600), .S(n601), .ZN(mantissa_ab_c[6]) );
  OAI21D4 U615 ( .A1(n557), .A2(n593), .B(n692), .ZN(mantissa_ab_c[17]) );
  CKMUX2D2 U616 ( .I0(c[14]), .I1(exp_ab[4]), .S(n897), .Z(exp_ab_c[4]) );
  MUX2ND2 U617 ( .I0(n617), .I1(n618), .S(n619), .ZN(mantissa_ab_c[2]) );
  OAI21D4 U618 ( .A1(n569), .A2(n593), .B(n728), .ZN(mantissa_ab_c[14]) );
  CKMUX2D2 U619 ( .I0(c[13]), .I1(exp_ab[3]), .S(n897), .Z(exp_ab_c[3]) );
  MUX2ND2 U620 ( .I0(n648), .I1(n649), .S(n650), .ZN(mantissa_ab_c[1]) );
  OAI21D4 U621 ( .A1(n577), .A2(n593), .B(n767), .ZN(mantissa_ab_c[11]) );
  MUX2ND2 U622 ( .I0(n898), .I1(n899), .S(n897), .ZN(exp_ab_c[2]) );
  OAI21D4 U623 ( .A1(n753), .A2(n593), .B(n754), .ZN(mantissa_ab_c[12]) );
  INVD1 U624 ( .I(fma_byp), .ZN(n593) );
  MUX2ND2 U625 ( .I0(n604), .I1(n605), .S(n606), .ZN(mantissa_ab_c[5]) );
  MUX2ND2 U626 ( .I0(n900), .I1(n901), .S(n897), .ZN(exp_ab_c[1]) );
  MUX2ND2 U627 ( .I0(n580), .I1(n581), .S(n582), .ZN(mantissa_ab_c[9]) );
  OA31D1 U628 ( .A1(n586), .A2(fma_byp), .A3(n584), .B(n587), .Z(n580) );
  MUX2ND2 U629 ( .I0(n902), .I1(n903), .S(n897), .ZN(exp_ab_c[0]) );
  MUX2ND2 U630 ( .I0(n608), .I1(n609), .S(n610), .ZN(mantissa_ab_c[4]) );
  OAI21D4 U631 ( .A1(n542), .A2(n543), .B(n544), .ZN(sign_ab_c) );
  OAI21D4 U632 ( .A1(n593), .A2(n576), .B(n778), .ZN(mantissa_ab_c[10]) );
  BUFFD2 U633 ( .I(n1147), .Z(mantissa_ab_c[21]) );
  ND2D1 U634 ( .A1(n585), .A2(n593), .ZN(n592) );
  NR2D3 U635 ( .A1(n651), .A2(fma_byp), .ZN(mantissa_ab_c[0]) );
  INVD1 U636 ( .I(n586), .ZN(n651) );
  TIEL U637 ( .ZN(n11) );
  MUX2ND0 U638 ( .I0(n545), .I1(c[15]), .S(fma_byp), .ZN(n544) );
  AOI31D0 U639 ( .A1(n546), .A2(n547), .A3(n548), .B(n549), .ZN(n545) );
  OAI21D0 U640 ( .A1(n550), .A2(n551), .B(n552), .ZN(n548) );
  CKND0 U641 ( .I(exp_ab_less), .ZN(n552) );
  OA31D0 U642 ( .A1(n551), .A2(exp_ab_greater), .A3(n550), .B(n553), .Z(n542)
         );
  NR2D0 U643 ( .A1(n554), .A2(c[9]), .ZN(n550) );
  AOI22D0 U644 ( .A1(n554), .A2(c[9]), .B1(n555), .B2(n556), .ZN(n551) );
  OAI221D0 U645 ( .A1(mantissa_ab[7]), .A2(n557), .B1(mantissa_ab[8]), .B2(
        n558), .C(n559), .ZN(n556) );
  OAI221D0 U646 ( .A1(c[6]), .A2(n560), .B1(c[7]), .B2(n561), .C(n562), .ZN(
        n559) );
  OAI221D0 U647 ( .A1(mantissa_ab[6]), .A2(n563), .B1(mantissa_ab[5]), .B2(
        n564), .C(n565), .ZN(n562) );
  OAI221D0 U648 ( .A1(c[4]), .A2(n566), .B1(c[5]), .B2(n567), .C(n568), .ZN(
        n565) );
  OAI222D0 U649 ( .A1(mantissa_ab[4]), .A2(n569), .B1(n570), .B2(n571), .C1(
        mantissa_ab[3]), .C2(n572), .ZN(n568) );
  MAOI222D0 U650 ( .A(n573), .B(n574), .C(c[2]), .ZN(n571) );
  AOI32D0 U651 ( .A1(n575), .A2(n576), .A3(mantissa_ab[0]), .B1(mantissa_ab[1]), .B2(n577), .ZN(n574) );
  CKND2D0 U652 ( .A1(c[1]), .A2(n578), .ZN(n575) );
  NR2D0 U653 ( .A1(c[3]), .A2(n579), .ZN(n570) );
  CKND2D0 U654 ( .A1(mantissa_ab[8]), .A2(n558), .ZN(n555) );
  AOI22D0 U655 ( .A1(n583), .A2(n584), .B1(mantissa_ab_c[0]), .B2(n585), .ZN(
        n581) );
  OR2D0 U656 ( .A1(n591), .A2(n592), .Z(n589) );
  AOI21D0 U657 ( .A1(n591), .A2(n593), .B(n594), .ZN(n588) );
  CKND2D0 U658 ( .A1(n583), .A2(n598), .ZN(n596) );
  CKND2D0 U659 ( .A1(n583), .A2(n602), .ZN(n600) );
  AOI21D0 U660 ( .A1(n603), .A2(n593), .B(n594), .ZN(n599) );
  OR2D0 U661 ( .A1(n607), .A2(n592), .Z(n605) );
  AOI21D0 U662 ( .A1(n607), .A2(n593), .B(n594), .ZN(n604) );
  AOI21D0 U663 ( .A1(n611), .A2(n593), .B(n594), .ZN(n609) );
  CKND2D0 U664 ( .A1(n583), .A2(n612), .ZN(n608) );
  IAO21D0 U665 ( .A1(n616), .A2(fma_byp), .B(n594), .ZN(n614) );
  CKND2D0 U666 ( .A1(n583), .A2(n620), .ZN(n618) );
  CKND0 U667 ( .I(n592), .ZN(n583) );
  AOI21D0 U668 ( .A1(n621), .A2(n593), .B(n594), .ZN(n617) );
  INR4D0 U669 ( .A1(n622), .B1(n623), .B2(n592), .B3(n624), .ZN(n1147) );
  CKND2D0 U670 ( .A1(n625), .A2(n626), .ZN(n623) );
  MUX2ND0 U671 ( .I0(n629), .I1(n630), .S(n624), .ZN(n628) );
  MUX2D0 U672 ( .I0(n631), .I1(n632), .S(n546), .Z(n624) );
  XNR2D0 U673 ( .A1(n633), .A2(n634), .ZN(n632) );
  AOI21D0 U674 ( .A1(n635), .A2(n636), .B(n637), .ZN(n633) );
  OAI21D0 U675 ( .A1(n638), .A2(n639), .B(n640), .ZN(n636) );
  AOI31D0 U676 ( .A1(n641), .A2(n642), .A3(n643), .B(n644), .ZN(n638) );
  CKND0 U677 ( .I(n645), .ZN(n635) );
  AO21D0 U678 ( .A1(n593), .A2(n646), .B(n594), .Z(n630) );
  NR2D0 U679 ( .A1(n646), .A2(n592), .ZN(n629) );
  INR2D0 U680 ( .A1(n625), .B1(n647), .ZN(n646) );
  CKND2D0 U681 ( .A1(mantissa_ab_c[0]), .A2(n585), .ZN(n649) );
  AOI21D0 U682 ( .A1(n651), .A2(n593), .B(n594), .ZN(n648) );
  MUX2ND0 U683 ( .I0(n654), .I1(n655), .S(n625), .ZN(n653) );
  MUX2ND0 U684 ( .I0(n656), .I1(n657), .S(add_byp), .ZN(n625) );
  CKXOR2D0 U685 ( .A1(n658), .A2(n645), .Z(n656) );
  AOI31D0 U686 ( .A1(n659), .A2(n660), .A3(n643), .B(n661), .ZN(n658) );
  OAI21D0 U687 ( .A1(n662), .A2(n663), .B(n664), .ZN(n660) );
  AOI21D0 U688 ( .A1(n665), .A2(n666), .B(n667), .ZN(n662) );
  INR2D0 U689 ( .A1(n647), .B1(n592), .ZN(n655) );
  OAI21D0 U690 ( .A1(fma_byp), .A2(n647), .B(n587), .ZN(n654) );
  ND4D0 U691 ( .A1(n622), .A2(n668), .A3(n669), .A4(n670), .ZN(n647) );
  MUX2ND0 U692 ( .I0(n672), .I1(n673), .S(n622), .ZN(n671) );
  MUX2ND0 U693 ( .I0(n674), .I1(n675), .S(add_byp), .ZN(n622) );
  CKXOR2D0 U694 ( .A1(n676), .A2(n639), .Z(n674) );
  AOI31D0 U695 ( .A1(n641), .A2(n677), .A3(n643), .B(n644), .ZN(n676) );
  OAI21D0 U696 ( .A1(n678), .A2(n664), .B(n679), .ZN(n644) );
  OAI21D0 U697 ( .A1(n680), .A2(n681), .B(n682), .ZN(n677) );
  CKND0 U698 ( .I(n683), .ZN(n681) );
  NR2D0 U699 ( .A1(n626), .A2(n592), .ZN(n673) );
  CKND0 U700 ( .I(n684), .ZN(n626) );
  OAI21D0 U701 ( .A1(fma_byp), .A2(n684), .B(n587), .ZN(n672) );
  CKND2D0 U702 ( .A1(n670), .A2(n685), .ZN(n684) );
  AN4D0 U703 ( .A1(n686), .A2(n687), .A3(n688), .A4(n689), .Z(n670) );
  AN2D0 U704 ( .A1(n690), .A2(n691), .Z(n689) );
  MUX2ND0 U705 ( .I0(n693), .I1(n694), .S(n687), .ZN(n692) );
  MUX2ND0 U706 ( .I0(n695), .I1(n696), .S(add_byp), .ZN(n687) );
  CKXOR2D0 U707 ( .A1(n697), .A2(n643), .Z(n695) );
  INR2D0 U708 ( .A1(n698), .B1(n592), .ZN(n694) );
  OAI21D0 U709 ( .A1(fma_byp), .A2(n698), .B(n587), .ZN(n693) );
  ND4D0 U710 ( .A1(n691), .A2(n688), .A3(n699), .A4(n700), .ZN(n698) );
  INR3D0 U711 ( .A1(n686), .B1(n584), .B2(n586), .ZN(n700) );
  ND4D0 U712 ( .A1(n619), .A2(n701), .A3(n702), .A4(n650), .ZN(n584) );
  NR2D0 U713 ( .A1(n615), .A2(n610), .ZN(n702) );
  MUX2ND0 U714 ( .I0(n704), .I1(n705), .S(n686), .ZN(n703) );
  MUX2ND0 U715 ( .I0(n706), .I1(n707), .S(add_byp), .ZN(n686) );
  CKXOR2D0 U716 ( .A1(n641), .A2(n642), .Z(n706) );
  CKND2D0 U717 ( .A1(n708), .A2(n682), .ZN(n642) );
  AOI32D0 U718 ( .A1(n665), .A2(n709), .A3(n710), .B1(n683), .B2(n711), .ZN(
        n708) );
  CKND0 U719 ( .I(n663), .ZN(n641) );
  NR2D0 U720 ( .A1(n712), .A2(n592), .ZN(n705) );
  AO21D0 U721 ( .A1(n593), .A2(n712), .B(n594), .Z(n704) );
  AN2D0 U722 ( .A1(n713), .A2(n691), .Z(n712) );
  MUX2ND0 U723 ( .I0(n715), .I1(n716), .S(n691), .ZN(n714) );
  MUX2ND0 U724 ( .I0(n717), .I1(n718), .S(add_byp), .ZN(n691) );
  CKXOR2D0 U725 ( .A1(n666), .A2(n665), .Z(n717) );
  OAI221D0 U726 ( .A1(n719), .A2(n720), .B1(n721), .B2(n722), .C(n723), .ZN(
        n666) );
  IND2D0 U727 ( .A1(n724), .B1(n725), .ZN(n722) );
  CKND0 U728 ( .I(n710), .ZN(n721) );
  NR2D0 U729 ( .A1(n726), .A2(n720), .ZN(n710) );
  NR2D0 U730 ( .A1(n713), .A2(n592), .ZN(n716) );
  IOA21D0 U731 ( .A1(n593), .A2(n713), .B(n587), .ZN(n715) );
  INR2D0 U732 ( .A1(n688), .B1(n727), .ZN(n713) );
  MUX2ND0 U733 ( .I0(n729), .I1(n730), .S(n688), .ZN(n728) );
  MUX2ND0 U734 ( .I0(n731), .I1(n732), .S(add_byp), .ZN(n688) );
  CKXOR2D0 U735 ( .A1(n680), .A2(n720), .Z(n731) );
  OA31D0 U736 ( .A1(n726), .A2(n733), .A3(n724), .B(n719), .Z(n680) );
  IAO21D0 U737 ( .A1(n726), .A2(n734), .B(n711), .ZN(n719) );
  OAI21D0 U738 ( .A1(n735), .A2(n736), .B(n737), .ZN(n711) );
  AOI21D0 U739 ( .A1(n738), .A2(n739), .B(n740), .ZN(n733) );
  OR2D0 U740 ( .A1(n735), .A2(n741), .Z(n726) );
  INR2D0 U741 ( .A1(n727), .B1(n592), .ZN(n730) );
  OAI21D0 U742 ( .A1(fma_byp), .A2(n727), .B(n587), .ZN(n729) );
  ND3D0 U743 ( .A1(n590), .A2(n591), .A3(n699), .ZN(n727) );
  AN3D0 U744 ( .A1(n690), .A2(n582), .A3(n742), .Z(n699) );
  INR2D0 U745 ( .A1(n597), .B1(n598), .ZN(n591) );
  CKND2D0 U746 ( .A1(n603), .A2(n601), .ZN(n598) );
  CKND0 U747 ( .I(n602), .ZN(n603) );
  CKND2D0 U748 ( .A1(n607), .A2(n606), .ZN(n602) );
  MUX2ND0 U749 ( .I0(n744), .I1(n745), .S(n690), .ZN(n743) );
  MUX2ND0 U750 ( .I0(n746), .I1(n747), .S(add_byp), .ZN(n690) );
  CKXOR2D0 U751 ( .A1(n735), .A2(n748), .Z(n746) );
  NR2D0 U752 ( .A1(n685), .A2(n592), .ZN(n745) );
  CKND0 U753 ( .I(n749), .ZN(n685) );
  OAI21D0 U754 ( .A1(fma_byp), .A2(n749), .B(n587), .ZN(n744) );
  CKND2D0 U755 ( .A1(n742), .A2(n750), .ZN(n749) );
  AN3D0 U756 ( .A1(n751), .A2(n752), .A3(n669), .Z(n742) );
  MUX2ND0 U757 ( .I0(n755), .I1(n756), .S(n669), .ZN(n754) );
  MUX2ND0 U758 ( .I0(n757), .I1(n758), .S(add_byp), .ZN(n669) );
  XNR2D0 U759 ( .A1(n741), .A2(n709), .ZN(n757) );
  OAI31D0 U760 ( .A1(n724), .A2(n759), .A3(n760), .B(n761), .ZN(n709) );
  CKND0 U761 ( .I(n762), .ZN(n761) );
  AOI21D0 U762 ( .A1(n763), .A2(n764), .B(n765), .ZN(n759) );
  NR2D0 U763 ( .A1(n668), .A2(n592), .ZN(n756) );
  AO21D0 U764 ( .A1(n593), .A2(n668), .B(n594), .Z(n755) );
  CKND0 U765 ( .I(n587), .ZN(n594) );
  INR2D0 U766 ( .A1(n752), .B1(n766), .ZN(n668) );
  MUX2ND0 U767 ( .I0(n768), .I1(n769), .S(n752), .ZN(n767) );
  MUX2ND0 U768 ( .I0(n770), .I1(n771), .S(add_byp), .ZN(n752) );
  XNR2D0 U769 ( .A1(n725), .A2(n724), .ZN(n770) );
  OAI21D0 U770 ( .A1(n772), .A2(n760), .B(n773), .ZN(n725) );
  CKND0 U771 ( .I(n738), .ZN(n760) );
  AOI21D0 U772 ( .A1(n774), .A2(n775), .B(n776), .ZN(n772) );
  CKND0 U773 ( .I(n777), .ZN(n776) );
  INR2D0 U774 ( .A1(n766), .B1(n592), .ZN(n769) );
  OAI21D0 U775 ( .A1(fma_byp), .A2(n766), .B(n587), .ZN(n768) );
  CKND2D0 U776 ( .A1(n750), .A2(n751), .ZN(n766) );
  MUX2ND0 U777 ( .I0(n779), .I1(n780), .S(n751), .ZN(n778) );
  MUX2ND0 U778 ( .I0(n781), .I1(n782), .S(add_byp), .ZN(n751) );
  CKXOR2D0 U779 ( .A1(n738), .A2(n739), .Z(n781) );
  OAI221D0 U780 ( .A1(n783), .A2(n784), .B1(n785), .B2(n786), .C(n777), .ZN(
        n739) );
  IAO21D0 U781 ( .A1(n787), .A2(n788), .B(n765), .ZN(n777) );
  NR2D0 U782 ( .A1(n789), .A2(n790), .ZN(n765) );
  CKND0 U783 ( .I(n774), .ZN(n784) );
  NR2D0 U784 ( .A1(n788), .A2(n791), .ZN(n774) );
  CKND0 U785 ( .I(n763), .ZN(n788) );
  NR2D0 U786 ( .A1(n790), .A2(n792), .ZN(n763) );
  AOI21D0 U787 ( .A1(n793), .A2(n794), .B(n795), .ZN(n783) );
  NR2D0 U788 ( .A1(n750), .A2(n592), .ZN(n780) );
  CKND0 U789 ( .I(n796), .ZN(n585) );
  CKND0 U790 ( .I(n797), .ZN(n750) );
  OAI21D0 U791 ( .A1(fma_byp), .A2(n797), .B(n587), .ZN(n779) );
  CKND2D0 U792 ( .A1(n796), .A2(n593), .ZN(n587) );
  XNR2D0 U793 ( .A1(n798), .A2(n799), .ZN(n796) );
  CKND2D0 U794 ( .A1(n800), .A2(n546), .ZN(n799) );
  CKXOR2D0 U795 ( .A1(n801), .A2(n802), .Z(n800) );
  AOI22D0 U796 ( .A1(n634), .A2(n803), .B1(n631), .B2(n804), .ZN(n801) );
  OAI21D0 U797 ( .A1(n805), .A2(n645), .B(n806), .ZN(n803) );
  CKND0 U798 ( .I(n637), .ZN(n806) );
  INR2D0 U799 ( .A1(n657), .B1(n807), .ZN(n637) );
  CKXOR2D0 U800 ( .A1(n807), .A2(n657), .Z(n645) );
  AOI31D0 U801 ( .A1(n659), .A2(n697), .A3(n643), .B(n661), .ZN(n805) );
  OAI21D0 U802 ( .A1(n639), .A2(n679), .B(n640), .ZN(n661) );
  CKND0 U803 ( .I(n678), .ZN(n643) );
  OAI21D0 U804 ( .A1(n696), .A2(n808), .B(n679), .ZN(n678) );
  CKND2D0 U805 ( .A1(n696), .A2(n808), .ZN(n679) );
  OAI21D0 U806 ( .A1(n809), .A2(n663), .B(n664), .ZN(n697) );
  OAI21D0 U807 ( .A1(n707), .A2(n810), .B(n664), .ZN(n663) );
  CKND2D0 U808 ( .A1(n707), .A2(n810), .ZN(n664) );
  AOI21D0 U809 ( .A1(n683), .A2(n811), .B(n812), .ZN(n809) );
  CKND0 U810 ( .I(n682), .ZN(n812) );
  IAO21D0 U811 ( .A1(n813), .A2(n723), .B(n667), .ZN(n682) );
  OAI21D0 U812 ( .A1(n748), .A2(n735), .B(n737), .ZN(n811) );
  OAI21D0 U813 ( .A1(n747), .A2(n814), .B(n737), .ZN(n735) );
  CKND2D0 U814 ( .A1(n747), .A2(n814), .ZN(n737) );
  OA21D0 U815 ( .A1(n815), .A2(n741), .B(n736), .Z(n748) );
  OAI21D0 U816 ( .A1(n758), .A2(n816), .B(n736), .ZN(n741) );
  CKND2D0 U817 ( .A1(n758), .A2(n816), .ZN(n736) );
  AOI31D0 U818 ( .A1(n738), .A2(n817), .A3(n818), .B(n762), .ZN(n815) );
  OAI21D0 U819 ( .A1(n773), .A2(n724), .B(n734), .ZN(n762) );
  AOI31D0 U820 ( .A1(n738), .A2(n819), .A3(n820), .B(n740), .ZN(n773) );
  NR2D0 U821 ( .A1(n724), .A2(n790), .ZN(n818) );
  OAI21D0 U822 ( .A1(n771), .A2(n821), .B(n734), .ZN(n724) );
  CKND2D0 U823 ( .A1(n771), .A2(n821), .ZN(n734) );
  CKND0 U824 ( .I(n822), .ZN(n821) );
  AOI21D0 U825 ( .A1(n823), .A2(n824), .B(n740), .ZN(n738) );
  NR2D0 U826 ( .A1(n823), .A2(n824), .ZN(n740) );
  NR2D0 U827 ( .A1(n720), .A2(n813), .ZN(n683) );
  CKND0 U828 ( .I(n665), .ZN(n813) );
  AOI21D0 U829 ( .A1(n825), .A2(n826), .B(n667), .ZN(n665) );
  NR2D0 U830 ( .A1(n825), .A2(n826), .ZN(n667) );
  OAI21D0 U831 ( .A1(n732), .A2(n827), .B(n723), .ZN(n720) );
  CKND2D0 U832 ( .A1(n732), .A2(n827), .ZN(n723) );
  CKND0 U833 ( .I(n828), .ZN(n827) );
  CKND0 U834 ( .I(n639), .ZN(n659) );
  OAI21D0 U835 ( .A1(n675), .A2(n829), .B(n640), .ZN(n639) );
  CKND2D0 U836 ( .A1(n675), .A2(n829), .ZN(n640) );
  CKXOR2D0 U837 ( .A1(n804), .A2(n631), .Z(n634) );
  ND3D0 U838 ( .A1(n582), .A2(n701), .A3(n607), .ZN(n797) );
  NR2D0 U839 ( .A1(n612), .A2(n610), .ZN(n607) );
  MUX2ND0 U840 ( .I0(n830), .I1(n831), .S(n546), .ZN(n610) );
  AO21D0 U841 ( .A1(n832), .A2(n833), .B(n834), .Z(n831) );
  CKND0 U842 ( .I(n611), .ZN(n612) );
  NR2D0 U843 ( .A1(n616), .A2(n615), .ZN(n611) );
  MUX2ND0 U844 ( .I0(n835), .I1(n836), .S(n546), .ZN(n615) );
  XNR2D0 U845 ( .A1(n837), .A2(n838), .ZN(n836) );
  CKND2D0 U846 ( .A1(n621), .A2(n619), .ZN(n616) );
  MUX2ND0 U847 ( .I0(n839), .I1(n840), .S(add_byp), .ZN(n619) );
  CKND0 U848 ( .I(n841), .ZN(n840) );
  CKXOR2D0 U849 ( .A1(n842), .A2(n843), .Z(n839) );
  CKND0 U850 ( .I(n620), .ZN(n621) );
  CKND2D0 U851 ( .A1(n650), .A2(n651), .ZN(n620) );
  CKXOR2D0 U852 ( .A1(n844), .A2(n845), .Z(n586) );
  CKXOR2D0 U853 ( .A1(n846), .A2(n847), .Z(n650) );
  CKND2D0 U854 ( .A1(n848), .A2(n546), .ZN(n847) );
  CKXOR2D0 U855 ( .A1(n849), .A2(n850), .Z(n848) );
  AN4D0 U856 ( .A1(n606), .A2(n601), .A3(n597), .A4(n590), .Z(n701) );
  MUX2ND0 U857 ( .I0(n851), .I1(n852), .S(add_byp), .ZN(n590) );
  XNR2D0 U858 ( .A1(n792), .A2(n764), .ZN(n851) );
  AO221D0 U859 ( .A1(n853), .A2(n854), .B1(n853), .B2(n834), .C(n855), .Z(n764) );
  MUX2ND0 U860 ( .I0(n856), .I1(n857), .S(add_byp), .ZN(n597) );
  XNR2D0 U861 ( .A1(n775), .A2(n791), .ZN(n856) );
  OAI31D0 U862 ( .A1(n858), .A2(n859), .A3(n860), .B(n861), .ZN(n775) );
  MUX2ND0 U863 ( .I0(n862), .I1(n863), .S(add_byp), .ZN(n601) );
  CKND0 U864 ( .I(n864), .ZN(n863) );
  CKXOR2D0 U865 ( .A1(n794), .A2(n793), .Z(n862) );
  OAI21D0 U866 ( .A1(n865), .A2(n860), .B(n866), .ZN(n794) );
  NR2D0 U867 ( .A1(n854), .A2(n834), .ZN(n865) );
  NR2D0 U868 ( .A1(n833), .A2(n832), .ZN(n834) );
  AOI21D0 U869 ( .A1(n867), .A2(n837), .B(n868), .ZN(n832) );
  OAI21D0 U870 ( .A1(n842), .A2(n843), .B(n869), .ZN(n867) );
  MAOI222D0 U871 ( .A(n846), .B(n870), .C(n850), .ZN(n843) );
  XNR2D0 U872 ( .A1(n871), .A2(n872), .ZN(n870) );
  CKND0 U873 ( .I(n873), .ZN(n842) );
  MUX2ND0 U874 ( .I0(n874), .I1(n875), .S(add_byp), .ZN(n606) );
  CKXOR2D0 U875 ( .A1(n860), .A2(n859), .Z(n874) );
  MUX2ND0 U876 ( .I0(n876), .I1(n820), .S(add_byp), .ZN(n582) );
  XNR2D0 U877 ( .A1(n790), .A2(n817), .ZN(n876) );
  OAI221D0 U878 ( .A1(n877), .A2(n792), .B1(n792), .B2(n878), .C(n789), .ZN(
        n817) );
  IND2D0 U879 ( .A1(n859), .B1(n853), .ZN(n878) );
  NR3D0 U880 ( .A1(n858), .A2(n860), .A3(n791), .ZN(n853) );
  OAI21D0 U881 ( .A1(n875), .A2(n879), .B(n866), .ZN(n860) );
  IAO21D0 U882 ( .A1(n880), .A2(n833), .B(n854), .ZN(n859) );
  AO21D0 U883 ( .A1(n830), .A2(n881), .B(n854), .Z(n833) );
  NR2D0 U884 ( .A1(n830), .A2(n881), .ZN(n854) );
  AOI21D0 U885 ( .A1(n837), .A2(n838), .B(n868), .ZN(n880) );
  OAI211D0 U886 ( .A1(n882), .A2(n883), .B(n884), .C(n869), .ZN(n838) );
  CKND0 U887 ( .I(n885), .ZN(n869) );
  OAI211D0 U888 ( .A1(n846), .A2(n849), .B(n873), .C(n850), .ZN(n884) );
  NR2D0 U889 ( .A1(n844), .A2(n886), .ZN(n850) );
  CKND0 U890 ( .I(n882), .ZN(n846) );
  CKND2D0 U891 ( .A1(n873), .A2(n849), .ZN(n883) );
  CKND0 U892 ( .I(n887), .ZN(n849) );
  AOI21D0 U893 ( .A1(n841), .A2(n888), .B(n885), .ZN(n873) );
  NR2D0 U894 ( .A1(n841), .A2(n888), .ZN(n885) );
  AOI21D0 U895 ( .A1(n835), .A2(n889), .B(n868), .ZN(n837) );
  NR2D0 U896 ( .A1(n835), .A2(n889), .ZN(n868) );
  IOA21D0 U897 ( .A1(n890), .A2(n891), .B(n789), .ZN(n792) );
  OR2D0 U898 ( .A1(n891), .A2(n890), .Z(n789) );
  CKND0 U899 ( .I(n852), .ZN(n890) );
  CKND0 U900 ( .I(n855), .ZN(n877) );
  OAI21D0 U901 ( .A1(n861), .A2(n791), .B(n787), .ZN(n855) );
  OAI21D0 U902 ( .A1(n857), .A2(n892), .B(n787), .ZN(n791) );
  CKND2D0 U903 ( .A1(n857), .A2(n892), .ZN(n787) );
  CKND0 U904 ( .I(n893), .ZN(n892) );
  CKND0 U905 ( .I(n894), .ZN(n857) );
  IAO21D0 U906 ( .A1(n858), .A2(n866), .B(n795), .ZN(n861) );
  CKND2D0 U907 ( .A1(n875), .A2(n879), .ZN(n866) );
  CKND0 U908 ( .I(n895), .ZN(n875) );
  CKND0 U909 ( .I(n793), .ZN(n858) );
  AOI21D0 U910 ( .A1(n864), .A2(n896), .B(n795), .ZN(n793) );
  NR2D0 U911 ( .A1(n864), .A2(n896), .ZN(n795) );
  XNR2D0 U912 ( .A1(n786), .A2(n785), .ZN(n790) );
  NR2D0 U913 ( .A1(fma_byp), .A2(n904), .ZN(n897) );
  NR2D0 U914 ( .A1(fma_byp), .A2(n785), .ZN(comp_mantissa_c[9]) );
  CKND0 U915 ( .I(n819), .ZN(n785) );
  CKXOR2D0 U916 ( .A1(n905), .A2(n906), .Z(n819) );
  NR2D0 U917 ( .A1(n907), .A2(n543), .ZN(n905) );
  NR2D0 U918 ( .A1(fma_byp), .A2(n891), .ZN(comp_mantissa_c[8]) );
  CKXOR2D0 U919 ( .A1(n908), .A2(n909), .Z(n891) );
  CKND2D0 U920 ( .A1(n910), .A2(n911), .ZN(n909) );
  NR2D0 U921 ( .A1(fma_byp), .A2(n893), .ZN(comp_mantissa_c[7]) );
  CKND2D0 U922 ( .A1(n912), .A2(n911), .ZN(n893) );
  MUX2ND0 U923 ( .I0(n543), .I1(n913), .S(n914), .ZN(n912) );
  AN2D0 U924 ( .A1(n915), .A2(n910), .Z(n913) );
  NR2D0 U925 ( .A1(fma_byp), .A2(n896), .ZN(comp_mantissa_c[6]) );
  CKND2D0 U926 ( .A1(n916), .A2(n915), .ZN(n896) );
  MUX2ND0 U927 ( .I0(n917), .I1(n543), .S(n918), .ZN(n916) );
  NR2D0 U928 ( .A1(n919), .A2(n543), .ZN(n917) );
  INR2D0 U929 ( .A1(n879), .B1(fma_byp), .ZN(comp_mantissa_c[5]) );
  INR2D0 U930 ( .A1(n920), .B1(n919), .ZN(n879) );
  MUX2ND0 U931 ( .I0(n921), .I1(n543), .S(n922), .ZN(n920) );
  NR2D0 U932 ( .A1(n923), .A2(n543), .ZN(n921) );
  NR2D0 U933 ( .A1(fma_byp), .A2(n881), .ZN(comp_mantissa_c[4]) );
  CKND2D0 U934 ( .A1(n924), .A2(n925), .ZN(n881) );
  MUX2ND0 U935 ( .I0(n926), .I1(n543), .S(n927), .ZN(n924) );
  NR2D0 U936 ( .A1(n928), .A2(n543), .ZN(n926) );
  NR2D0 U937 ( .A1(fma_byp), .A2(n889), .ZN(comp_mantissa_c[3]) );
  CKND2D0 U938 ( .A1(n929), .A2(n930), .ZN(n889) );
  MUX2ND0 U939 ( .I0(n931), .I1(n543), .S(n932), .ZN(n929) );
  NR2D0 U940 ( .A1(n933), .A2(n543), .ZN(n931) );
  NR2D0 U941 ( .A1(fma_byp), .A2(n888), .ZN(comp_mantissa_c[2]) );
  CKND2D0 U942 ( .A1(n934), .A2(n935), .ZN(n888) );
  MUX2ND0 U943 ( .I0(n936), .I1(n543), .S(n937), .ZN(n934) );
  OAI22D0 U944 ( .A1(n938), .A2(n845), .B1(n543), .B2(n871), .ZN(n936) );
  NR2D0 U945 ( .A1(fma_byp), .A2(n802), .ZN(comp_mantissa_c[21]) );
  OAI31D0 U946 ( .A1(n939), .A2(n940), .A3(n941), .B(n910), .ZN(n802) );
  ND3D0 U947 ( .A1(n942), .A2(n943), .A3(n944), .ZN(n939) );
  MUX2D0 U948 ( .I0(n945), .I1(n804), .S(n593), .Z(comp_mantissa_c[20]) );
  XNR2D0 U949 ( .A1(n946), .A2(n944), .ZN(n804) );
  OAI211D0 U950 ( .A1(n947), .A2(n547), .B(n948), .C(n945), .ZN(n944) );
  AOI21D0 U951 ( .A1(n949), .A2(n950), .B(n938), .ZN(n946) );
  OR2D0 U952 ( .A1(n942), .A2(add_byp), .Z(n950) );
  NR2D0 U953 ( .A1(fma_byp), .A2(n887), .ZN(comp_mantissa_c[1]) );
  CKXOR2D0 U954 ( .A1(n872), .A2(n871), .Z(n887) );
  NR2D0 U955 ( .A1(n938), .A2(n845), .ZN(n872) );
  OR2D0 U956 ( .A1(n886), .A2(add_byp), .Z(n845) );
  MUX2ND0 U957 ( .I0(n807), .I1(n652), .S(fma_byp), .ZN(comp_mantissa_c[19])
         );
  CKXOR2D0 U958 ( .A1(n951), .A2(n942), .Z(n807) );
  CKND2D0 U959 ( .A1(n952), .A2(n948), .ZN(n942) );
  MUX2ND0 U960 ( .I0(n652), .I1(n953), .S(exp_ab_greater), .ZN(n952) );
  NR2D0 U961 ( .A1(n938), .A2(n949), .ZN(n951) );
  OAI31D0 U962 ( .A1(n954), .A2(n940), .A3(n955), .B(n546), .ZN(n949) );
  CKND2D0 U963 ( .A1(n956), .A2(n943), .ZN(n954) );
  CKND0 U964 ( .I(c[15]), .ZN(n938) );
  MUX2D0 U965 ( .I0(c[8]), .I1(n829), .S(n593), .Z(comp_mantissa_c[18]) );
  XNR2D0 U966 ( .A1(n957), .A2(n943), .ZN(n829) );
  CKND2D0 U967 ( .A1(n958), .A2(n948), .ZN(n943) );
  MUX2ND0 U968 ( .I0(n558), .I1(n959), .S(exp_ab_greater), .ZN(n958) );
  IAO21D0 U969 ( .A1(n941), .A2(n940), .B(n543), .ZN(n957) );
  CKND2D0 U970 ( .A1(n960), .A2(n961), .ZN(n940) );
  MUX2D0 U971 ( .I0(c[7]), .I1(n808), .S(n593), .Z(comp_mantissa_c[17]) );
  XNR2D0 U972 ( .A1(n962), .A2(n961), .ZN(n808) );
  CKND2D0 U973 ( .A1(n963), .A2(n948), .ZN(n961) );
  CKND2D0 U974 ( .A1(exp_ab_greater), .A2(n964), .ZN(n948) );
  MUX2ND0 U975 ( .I0(n557), .I1(n965), .S(exp_ab_greater), .ZN(n963) );
  AOI31D0 U976 ( .A1(n907), .A2(n960), .A3(n966), .B(n543), .ZN(n962) );
  NR2D0 U977 ( .A1(n906), .A2(n967), .ZN(n966) );
  IINR4D0 U978 ( .A1(n968), .A2(n969), .B1(n970), .B2(n971), .ZN(n960) );
  NR2D0 U979 ( .A1(n911), .A2(n908), .ZN(n907) );
  IND2D0 U980 ( .A1(n915), .B1(n972), .ZN(n911) );
  CKND2D0 U981 ( .A1(n919), .A2(n918), .ZN(n915) );
  AN2D0 U982 ( .A1(n922), .A2(n923), .Z(n919) );
  MUX2D0 U983 ( .I0(c[6]), .I1(n810), .S(n593), .Z(comp_mantissa_c[16]) );
  CKXOR2D0 U984 ( .A1(n973), .A2(n970), .Z(n810) );
  MUX2ND0 U985 ( .I0(n563), .I1(n974), .S(exp_ab_greater), .ZN(n970) );
  CKND2D0 U986 ( .A1(n975), .A2(n976), .ZN(n974) );
  INR2D0 U987 ( .A1(n977), .B1(n543), .ZN(n973) );
  MUX2ND0 U988 ( .I0(n826), .I1(n564), .S(fma_byp), .ZN(comp_mantissa_c[15])
         );
  CKND2D0 U989 ( .A1(n978), .A2(n977), .ZN(n826) );
  CKND2D0 U990 ( .A1(n979), .A2(n969), .ZN(n977) );
  MUX2ND0 U991 ( .I0(n969), .I1(n980), .S(n910), .ZN(n978) );
  NR2D0 U992 ( .A1(n979), .A2(n969), .ZN(n980) );
  CKND0 U993 ( .I(n981), .ZN(n979) );
  MUX2D0 U994 ( .I0(n982), .I1(n564), .S(n547), .Z(n969) );
  AOI22D0 U995 ( .A1(n983), .A2(n984), .B1(n985), .B2(n986), .ZN(n982) );
  MUX2ND0 U996 ( .I0(n828), .I1(n569), .S(fma_byp), .ZN(comp_mantissa_c[14])
         );
  CKND2D0 U997 ( .A1(n987), .A2(n981), .ZN(n828) );
  CKND2D0 U998 ( .A1(n988), .A2(n968), .ZN(n981) );
  MUX2ND0 U999 ( .I0(n968), .I1(n989), .S(n910), .ZN(n987) );
  NR2D0 U1000 ( .A1(n988), .A2(n968), .ZN(n989) );
  NR2D0 U1001 ( .A1(n941), .A2(n971), .ZN(n988) );
  MUX2D0 U1002 ( .I0(n990), .I1(n569), .S(n547), .Z(n968) );
  AOI22D0 U1003 ( .A1(n983), .A2(n991), .B1(n985), .B2(n992), .ZN(n990) );
  MUX2D0 U1004 ( .I0(c[3]), .I1(n814), .S(n593), .Z(comp_mantissa_c[13]) );
  CKXOR2D0 U1005 ( .A1(n993), .A2(n971), .Z(n814) );
  MUX2ND0 U1006 ( .I0(n572), .I1(n994), .S(exp_ab_greater), .ZN(n971) );
  AOI22D0 U1007 ( .A1(n983), .A2(n995), .B1(n985), .B2(n996), .ZN(n994) );
  AN2D0 U1008 ( .A1(n941), .A2(n910), .Z(n993) );
  IND2D0 U1009 ( .A1(n967), .B1(n997), .ZN(n941) );
  ND3D0 U1010 ( .A1(n956), .A2(n998), .A3(n999), .ZN(n967) );
  MUX2D0 U1011 ( .I0(c[2]), .I1(n816), .S(n593), .Z(comp_mantissa_c[12]) );
  XNR2D0 U1012 ( .A1(n1000), .A2(n956), .ZN(n816) );
  MUX2D0 U1013 ( .I0(n1001), .I1(n753), .S(n547), .Z(n956) );
  AOI222D0 U1014 ( .A1(n947), .A2(n1002), .B1(n985), .B2(n1003), .C1(n983), 
        .C2(n1004), .ZN(n1001) );
  INR2D0 U1015 ( .A1(n955), .B1(n543), .ZN(n1000) );
  MUX2ND0 U1016 ( .I0(n822), .I1(n577), .S(fma_byp), .ZN(comp_mantissa_c[11])
         );
  CKND2D0 U1017 ( .A1(n1005), .A2(n955), .ZN(n822) );
  CKND2D0 U1018 ( .A1(n1006), .A2(n999), .ZN(n955) );
  MUX2ND0 U1019 ( .I0(n999), .I1(n1007), .S(n910), .ZN(n1005) );
  NR2D0 U1020 ( .A1(n1006), .A2(n999), .ZN(n1007) );
  CKND0 U1021 ( .I(n1008), .ZN(n1006) );
  MUX2D0 U1022 ( .I0(n1009), .I1(n577), .S(n547), .Z(n999) );
  AOI222D0 U1023 ( .A1(n983), .A2(n986), .B1(n1002), .B2(n984), .C1(n985), 
        .C2(n1010), .ZN(n1009) );
  MUX2ND0 U1024 ( .I0(n824), .I1(n576), .S(fma_byp), .ZN(comp_mantissa_c[10])
         );
  CKND2D0 U1025 ( .A1(n1011), .A2(n1008), .ZN(n824) );
  CKND2D0 U1026 ( .A1(n997), .A2(n998), .ZN(n1008) );
  MUX2ND0 U1027 ( .I0(n998), .I1(n1012), .S(n910), .ZN(n1011) );
  CKND0 U1028 ( .I(n543), .ZN(n910) );
  CKND2D0 U1029 ( .A1(c[15]), .A2(n546), .ZN(n543) );
  CKND0 U1030 ( .I(add_byp), .ZN(n546) );
  NR2D0 U1031 ( .A1(n997), .A2(n998), .ZN(n1012) );
  AN4D0 U1032 ( .A1(n922), .A2(n918), .A3(n923), .A4(n1013), .Z(n997) );
  NR3D0 U1033 ( .A1(n914), .A2(n906), .A3(n908), .ZN(n1013) );
  AN2D0 U1034 ( .A1(n1014), .A2(exp_ab_greater), .Z(n908) );
  OAI222D0 U1035 ( .A1(n1015), .A2(n964), .B1(n1016), .B2(n1017), .C1(n1018), 
        .C2(n1019), .ZN(n1014) );
  CKND2D0 U1036 ( .A1(n976), .A2(n1020), .ZN(n1017) );
  AN2D0 U1037 ( .A1(n1021), .A2(exp_ab_greater), .Z(n906) );
  OAI222D0 U1038 ( .A1(n965), .A2(n1022), .B1(n1023), .B2(n964), .C1(n1024), 
        .C2(n1019), .ZN(n1021) );
  CKND0 U1039 ( .I(n972), .ZN(n914) );
  CKND2D0 U1040 ( .A1(exp_ab_greater), .A2(n1025), .ZN(n972) );
  OAI221D0 U1041 ( .A1(n1026), .A2(n1019), .B1(n1027), .B2(n1022), .C(n1028), 
        .ZN(n1025) );
  OA32D0 U1042 ( .A1(n576), .A2(n1029), .A3(n964), .B1(n1030), .B2(n953), .Z(
        n1028) );
  CKND0 U1043 ( .I(n925), .ZN(n923) );
  CKND2D0 U1044 ( .A1(n928), .A2(n927), .ZN(n925) );
  CKND2D0 U1045 ( .A1(exp_ab_greater), .A2(n1031), .ZN(n927) );
  OAI221D0 U1046 ( .A1(n1018), .A2(n1022), .B1(n1032), .B2(n1030), .C(n1033), 
        .ZN(n1031) );
  MAOI22D0 U1047 ( .A1(n947), .A2(n1034), .B1(n1019), .B2(n1015), .ZN(n1033)
         );
  CKND0 U1048 ( .I(n1004), .ZN(n1032) );
  CKND0 U1049 ( .I(n930), .ZN(n928) );
  CKND2D0 U1050 ( .A1(n933), .A2(n932), .ZN(n930) );
  CKND2D0 U1051 ( .A1(exp_ab_greater), .A2(n1035), .ZN(n932) );
  OAI221D0 U1052 ( .A1(n1026), .A2(n1022), .B1(n1027), .B2(n1030), .C(n1036), 
        .ZN(n1035) );
  AOI32D0 U1053 ( .A1(c[0]), .A2(n1037), .A3(n983), .B1(n1034), .B2(n984), 
        .ZN(n1036) );
  CKND0 U1054 ( .I(n953), .ZN(n984) );
  AOI22D0 U1055 ( .A1(c[9]), .A2(n1038), .B1(n945), .B2(n1039), .ZN(n953) );
  CKND0 U1056 ( .I(n1040), .ZN(n1034) );
  CKND0 U1057 ( .I(n986), .ZN(n1027) );
  OAI221D0 U1058 ( .A1(n558), .A2(n1029), .B1(n564), .B2(n1041), .C(n1042), 
        .ZN(n986) );
  AOI22D0 U1059 ( .A1(n1043), .A2(c[7]), .B1(n1039), .B2(c[6]), .ZN(n1042) );
  CKND0 U1060 ( .I(c[8]), .ZN(n558) );
  CKND0 U1061 ( .I(n1010), .ZN(n1026) );
  OAI221D0 U1062 ( .A1(n569), .A2(n1029), .B1(n577), .B2(n1041), .C(n1044), 
        .ZN(n1010) );
  AOI22D0 U1063 ( .A1(n1043), .A2(c[3]), .B1(n1039), .B2(c[2]), .ZN(n1044) );
  CKND0 U1064 ( .I(c[1]), .ZN(n577) );
  CKND0 U1065 ( .I(n935), .ZN(n933) );
  ND3D0 U1066 ( .A1(n937), .A2(n886), .A3(n871), .ZN(n935) );
  CKND2D0 U1067 ( .A1(exp_ab_greater), .A2(n1045), .ZN(n871) );
  OAI222D0 U1068 ( .A1(n965), .A2(n1040), .B1(n1023), .B2(n1022), .C1(n1024), 
        .C2(n1030), .ZN(n1045) );
  CKND2D0 U1069 ( .A1(exp_ab_greater), .A2(n1046), .ZN(n937) );
  OAI222D0 U1070 ( .A1(n1047), .A2(n1022), .B1(n959), .B2(n1040), .C1(n1048), 
        .C2(n1030), .ZN(n1046) );
  ND3D0 U1071 ( .A1(n1049), .A2(n1016), .A3(exp_diff[4]), .ZN(n1040) );
  CKND2D0 U1072 ( .A1(exp_ab_greater), .A2(n1050), .ZN(n918) );
  OAI222D0 U1073 ( .A1(n1047), .A2(n1019), .B1(n959), .B2(n1030), .C1(n1048), 
        .C2(n1022), .ZN(n1050) );
  CKND0 U1074 ( .I(n992), .ZN(n1048) );
  CKND0 U1075 ( .I(n1051), .ZN(n1047) );
  CKND2D0 U1076 ( .A1(exp_ab_greater), .A2(n1052), .ZN(n922) );
  OAI222D0 U1077 ( .A1(n965), .A2(n1030), .B1(n1023), .B2(n1019), .C1(n1024), 
        .C2(n1022), .ZN(n1052) );
  CKND0 U1078 ( .I(n996), .ZN(n1024) );
  OAI221D0 U1079 ( .A1(n563), .A2(n1029), .B1(n572), .B2(n1041), .C(n1053), 
        .ZN(n996) );
  AOI22D0 U1080 ( .A1(n1043), .A2(c[5]), .B1(n1039), .B2(c[4]), .ZN(n1053) );
  AOI222D0 U1081 ( .A1(n1039), .A2(c[0]), .B1(c[1]), .B2(n1043), .C1(c[2]), 
        .C2(n1037), .ZN(n1023) );
  CKND0 U1082 ( .I(n995), .ZN(n965) );
  OAI221D0 U1083 ( .A1(n557), .A2(n1041), .B1(n627), .B2(n1029), .C(n1054), 
        .ZN(n995) );
  AOI22D0 U1084 ( .A1(n1043), .A2(c[9]), .B1(n1039), .B2(c[8]), .ZN(n1054) );
  MUX2D0 U1085 ( .I0(n1055), .I1(n576), .S(n547), .Z(n998) );
  AOI222D0 U1086 ( .A1(n983), .A2(n992), .B1(n1002), .B2(n991), .C1(n985), 
        .C2(n1051), .ZN(n1055) );
  OAI221D0 U1087 ( .A1(n572), .A2(n1029), .B1(n1041), .B2(n576), .C(n1056), 
        .ZN(n1051) );
  AOI22D0 U1088 ( .A1(n1043), .A2(c[2]), .B1(n1039), .B2(c[1]), .ZN(n1056) );
  CKND0 U1089 ( .I(c[0]), .ZN(n576) );
  CKND0 U1090 ( .I(c[3]), .ZN(n572) );
  CKND0 U1091 ( .I(n964), .ZN(n985) );
  CKND2D0 U1092 ( .A1(n975), .A2(n1049), .ZN(n964) );
  CKND0 U1093 ( .I(n959), .ZN(n991) );
  AOI222D0 U1094 ( .A1(c[8]), .A2(n1038), .B1(c[9]), .B2(n1039), .C1(n945), 
        .C2(n1043), .ZN(n959) );
  CKND0 U1095 ( .I(n1022), .ZN(n1002) );
  OAI221D0 U1096 ( .A1(n557), .A2(n1029), .B1(n569), .B2(n1041), .C(n1057), 
        .ZN(n992) );
  AOI22D0 U1097 ( .A1(n1043), .A2(c[6]), .B1(n1039), .B2(c[5]), .ZN(n1057) );
  CKND0 U1098 ( .I(c[4]), .ZN(n569) );
  CKND0 U1099 ( .I(c[7]), .ZN(n557) );
  CKND0 U1100 ( .I(n1019), .ZN(n983) );
  CKND2D0 U1101 ( .A1(n975), .A2(exp_diff[2]), .ZN(n1019) );
  NR2D0 U1102 ( .A1(exp_diff[4]), .A2(exp_diff[3]), .ZN(n975) );
  NR2D0 U1103 ( .A1(fma_byp), .A2(n886), .ZN(comp_mantissa_c[0]) );
  CKND2D0 U1104 ( .A1(exp_ab_greater), .A2(n1058), .ZN(n886) );
  OAI222D0 U1105 ( .A1(n1015), .A2(n1022), .B1(n1020), .B2(n1059), .C1(n1018), 
        .C2(n1030), .ZN(n1058) );
  ND3D0 U1106 ( .A1(exp_diff[2]), .A2(n1020), .A3(exp_diff[3]), .ZN(n1030) );
  CKND0 U1107 ( .I(n1003), .ZN(n1018) );
  OAI221D0 U1108 ( .A1(n564), .A2(n1029), .B1(n753), .B2(n1041), .C(n1060), 
        .ZN(n1003) );
  AOI22D0 U1109 ( .A1(n1043), .A2(c[4]), .B1(n1039), .B2(c[3]), .ZN(n1060) );
  CKND0 U1110 ( .I(c[2]), .ZN(n753) );
  CKND0 U1111 ( .I(c[5]), .ZN(n564) );
  CKND2D0 U1112 ( .A1(n976), .A2(n1016), .ZN(n1059) );
  CKND0 U1113 ( .I(exp_diff[3]), .ZN(n1016) );
  MUX2D0 U1114 ( .I0(n947), .I1(n1004), .S(n1049), .Z(n976) );
  OAI221D0 U1115 ( .A1(n652), .A2(n1029), .B1(n563), .B2(n1041), .C(n1061), 
        .ZN(n1004) );
  AOI22D0 U1116 ( .A1(n1043), .A2(c[8]), .B1(n1039), .B2(c[7]), .ZN(n1061) );
  INR2D0 U1117 ( .A1(exp_diff[0]), .B1(exp_diff[1]), .ZN(n1039) );
  CKND0 U1118 ( .I(c[6]), .ZN(n563) );
  CKND0 U1119 ( .I(c[9]), .ZN(n652) );
  NR2D0 U1120 ( .A1(n1041), .A2(n627), .ZN(n947) );
  CKND0 U1121 ( .I(n945), .ZN(n627) );
  ND4D0 U1122 ( .A1(n902), .A2(n900), .A3(n1062), .A4(n898), .ZN(n945) );
  CKND0 U1123 ( .I(c[12]), .ZN(n898) );
  NR2D0 U1124 ( .A1(c[14]), .A2(c[13]), .ZN(n1062) );
  CKND0 U1125 ( .I(c[11]), .ZN(n900) );
  CKND0 U1126 ( .I(c[10]), .ZN(n902) );
  CKND0 U1127 ( .I(n1038), .ZN(n1041) );
  NR2D0 U1128 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n1038) );
  ND3D0 U1129 ( .A1(n1049), .A2(n1020), .A3(exp_diff[3]), .ZN(n1022) );
  CKND0 U1130 ( .I(exp_diff[4]), .ZN(n1020) );
  CKND0 U1131 ( .I(exp_diff[2]), .ZN(n1049) );
  AOI22D0 U1132 ( .A1(c[1]), .A2(n1037), .B1(n1043), .B2(c[0]), .ZN(n1015) );
  INR2D0 U1133 ( .A1(exp_diff[1]), .B1(exp_diff[0]), .ZN(n1043) );
  CKND0 U1134 ( .I(n1029), .ZN(n1037) );
  CKND2D0 U1135 ( .A1(exp_diff[0]), .A2(exp_diff[1]), .ZN(n1029) );
  MUX2ND0 U1136 ( .I0(n786), .I1(n554), .S(fma_byp), .ZN(comp_mantissa_ab[9])
         );
  CKND0 U1137 ( .I(mantissa_ab[9]), .ZN(n554) );
  CKND0 U1138 ( .I(n820), .ZN(n786) );
  XNR2D0 U1139 ( .A1(n1063), .A2(n1064), .ZN(n820) );
  NR2D0 U1140 ( .A1(n1065), .A2(n549), .ZN(n1063) );
  MUX2D0 U1141 ( .I0(mantissa_ab[8]), .I1(n852), .S(n593), .Z(
        comp_mantissa_ab[8]) );
  XNR2D0 U1142 ( .A1(n1066), .A2(n1067), .ZN(n852) );
  NR2D0 U1143 ( .A1(n1068), .A2(n549), .ZN(n1066) );
  MUX2ND0 U1144 ( .I0(n894), .I1(n561), .S(fma_byp), .ZN(comp_mantissa_ab[7])
         );
  CKND0 U1145 ( .I(mantissa_ab[7]), .ZN(n561) );
  CKND2D0 U1146 ( .A1(n1069), .A2(n1070), .ZN(n894) );
  MUX2ND0 U1147 ( .I0(n1071), .I1(n1072), .S(sign_ab), .ZN(n1069) );
  NR2D0 U1148 ( .A1(n1073), .A2(n1071), .ZN(n1072) );
  MUX2ND0 U1149 ( .I0(n864), .I1(n560), .S(fma_byp), .ZN(comp_mantissa_ab[6])
         );
  CKND0 U1150 ( .I(mantissa_ab[6]), .ZN(n560) );
  CKND2D0 U1151 ( .A1(n1074), .A2(n1075), .ZN(n864) );
  MUX2ND0 U1152 ( .I0(n1076), .I1(n1077), .S(sign_ab), .ZN(n1074) );
  NR2D0 U1153 ( .A1(n1078), .A2(n1076), .ZN(n1077) );
  MUX2ND0 U1154 ( .I0(n895), .I1(n567), .S(fma_byp), .ZN(comp_mantissa_ab[5])
         );
  CKND0 U1155 ( .I(mantissa_ab[5]), .ZN(n567) );
  CKND2D0 U1156 ( .A1(n1079), .A2(n1080), .ZN(n895) );
  MUX2ND0 U1157 ( .I0(n1081), .I1(n1082), .S(sign_ab), .ZN(n1079) );
  NR2D0 U1158 ( .A1(n1083), .A2(n1081), .ZN(n1082) );
  MUX2ND0 U1159 ( .I0(n830), .I1(n566), .S(fma_byp), .ZN(comp_mantissa_ab[4])
         );
  CKND0 U1160 ( .I(mantissa_ab[4]), .ZN(n566) );
  CKND2D0 U1161 ( .A1(n1084), .A2(n1085), .ZN(n830) );
  MUX2ND0 U1162 ( .I0(n1086), .I1(n1087), .S(sign_ab), .ZN(n1084) );
  NR2D0 U1163 ( .A1(n1088), .A2(n1086), .ZN(n1087) );
  MUX2ND0 U1164 ( .I0(n835), .I1(n579), .S(fma_byp), .ZN(comp_mantissa_ab[3])
         );
  CKND0 U1165 ( .I(mantissa_ab[3]), .ZN(n579) );
  CKND2D0 U1166 ( .A1(n1089), .A2(n1090), .ZN(n835) );
  MUX2ND0 U1167 ( .I0(n1091), .I1(n1092), .S(sign_ab), .ZN(n1089) );
  NR2D0 U1168 ( .A1(n1093), .A2(n1091), .ZN(n1092) );
  MUX2ND0 U1169 ( .I0(n841), .I1(n573), .S(fma_byp), .ZN(comp_mantissa_ab[2])
         );
  CKND0 U1170 ( .I(mantissa_ab[2]), .ZN(n573) );
  IND2D0 U1171 ( .A1(n1093), .B1(n1094), .ZN(n841) );
  MUX2ND0 U1172 ( .I0(n1095), .I1(n1096), .S(sign_ab), .ZN(n1094) );
  INR2D0 U1173 ( .A1(n1097), .B1(n1095), .ZN(n1096) );
  NR2D0 U1174 ( .A1(fma_byp), .A2(n798), .ZN(comp_mantissa_ab[21]) );
  OAI31D0 U1175 ( .A1(n1098), .A2(n1099), .A3(n1100), .B(sign_ab), .ZN(n798)
         );
  CKND2D0 U1176 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
  MUX2D0 U1177 ( .I0(N800), .I1(n631), .S(n593), .Z(comp_mantissa_ab[20]) );
  CKXOR2D0 U1178 ( .A1(n1103), .A2(n1099), .Z(n631) );
  MUX2D0 U1179 ( .I0(N800), .I1(N65), .S(n904), .Z(n1099) );
  AOI21D0 U1180 ( .A1(n1104), .A2(n1101), .B(n549), .ZN(n1103) );
  MUX2ND0 U1181 ( .I0(n882), .I1(n578), .S(fma_byp), .ZN(comp_mantissa_ab[1])
         );
  CKND0 U1182 ( .I(mantissa_ab[1]), .ZN(n578) );
  CKND2D0 U1183 ( .A1(n1105), .A2(n1097), .ZN(n882) );
  MUX2ND0 U1184 ( .I0(n1106), .I1(n1107), .S(sign_ab), .ZN(n1105) );
  NR2D0 U1185 ( .A1(n844), .A2(n1106), .ZN(n1107) );
  MUX2D0 U1186 ( .I0(mantissa_ab[19]), .I1(n657), .S(n593), .Z(
        comp_mantissa_ab[19]) );
  XNR2D0 U1187 ( .A1(n1108), .A2(n1101), .ZN(n657) );
  MUX2ND0 U1188 ( .I0(mantissa_ab[19]), .I1(N64), .S(n904), .ZN(n1101) );
  NR2D0 U1189 ( .A1(n1104), .A2(n549), .ZN(n1108) );
  AN4D0 U1190 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1102), .Z(n1104) );
  MUX2D0 U1191 ( .I0(mantissa_ab[18]), .I1(n675), .S(n593), .Z(
        comp_mantissa_ab[18]) );
  XNR2D0 U1192 ( .A1(n1112), .A2(n1102), .ZN(n675) );
  MUX2ND0 U1193 ( .I0(mantissa_ab[18]), .I1(N63), .S(n904), .ZN(n1102) );
  INR2D0 U1194 ( .A1(n1100), .B1(n549), .ZN(n1112) );
  CKND2D0 U1195 ( .A1(n1110), .A2(n1113), .ZN(n1100) );
  INR2D0 U1196 ( .A1(n1114), .B1(n1115), .ZN(n1110) );
  MUX2D0 U1197 ( .I0(mantissa_ab[17]), .I1(n696), .S(n593), .Z(
        comp_mantissa_ab[17]) );
  XNR2D0 U1198 ( .A1(n1116), .A2(n1114), .ZN(n696) );
  MUX2ND0 U1199 ( .I0(mantissa_ab[17]), .I1(N62), .S(n904), .ZN(n1114) );
  AOI31D0 U1200 ( .A1(n1065), .A2(n1117), .A3(n1118), .B(n549), .ZN(n1116) );
  INR2D0 U1201 ( .A1(n1064), .B1(n1115), .ZN(n1118) );
  ND4D0 U1202 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1115) );
  AN4D0 U1203 ( .A1(n1086), .A2(n1091), .A3(n1123), .A4(n1124), .Z(n1065) );
  AN3D0 U1204 ( .A1(n1095), .A2(n844), .A3(n1106), .Z(n1124) );
  MUX2D0 U1205 ( .I0(mantissa_ab[16]), .I1(n707), .S(n593), .Z(
        comp_mantissa_ab[16]) );
  XNR2D0 U1206 ( .A1(n1125), .A2(n1119), .ZN(n707) );
  MUX2ND0 U1207 ( .I0(mantissa_ab[16]), .I1(N61), .S(n904), .ZN(n1119) );
  INR2D0 U1208 ( .A1(n1126), .B1(n549), .ZN(n1125) );
  MUX2D0 U1209 ( .I0(mantissa_ab[15]), .I1(n718), .S(n593), .Z(
        comp_mantissa_ab[15]) );
  CKND0 U1210 ( .I(n825), .ZN(n718) );
  CKND2D0 U1211 ( .A1(n1127), .A2(n1126), .ZN(n825) );
  CKND2D0 U1212 ( .A1(n1128), .A2(n1120), .ZN(n1126) );
  MUX2ND0 U1213 ( .I0(n1120), .I1(n1129), .S(sign_ab), .ZN(n1127) );
  NR2D0 U1214 ( .A1(n1128), .A2(n1120), .ZN(n1129) );
  MUX2ND0 U1215 ( .I0(N60), .I1(mantissa_ab[15]), .S(n553), .ZN(n1120) );
  MUX2D0 U1216 ( .I0(mantissa_ab[14]), .I1(n732), .S(n593), .Z(
        comp_mantissa_ab[14]) );
  INR2D0 U1217 ( .A1(n1130), .B1(n1128), .ZN(n732) );
  AN2D0 U1218 ( .A1(n1131), .A2(n1121), .Z(n1128) );
  MUX2ND0 U1219 ( .I0(n1121), .I1(n1132), .S(sign_ab), .ZN(n1130) );
  NR2D0 U1220 ( .A1(n1131), .A2(n1121), .ZN(n1132) );
  AN4D0 U1221 ( .A1(n1068), .A2(n1117), .A3(n1133), .A4(n1064), .Z(n1131) );
  AN2D0 U1222 ( .A1(n1067), .A2(n1122), .Z(n1133) );
  CKND0 U1223 ( .I(n1070), .ZN(n1068) );
  CKND2D0 U1224 ( .A1(n1073), .A2(n1071), .ZN(n1070) );
  CKND0 U1225 ( .I(n1075), .ZN(n1073) );
  CKND2D0 U1226 ( .A1(n1078), .A2(n1076), .ZN(n1075) );
  CKND0 U1227 ( .I(n1080), .ZN(n1078) );
  CKND2D0 U1228 ( .A1(n1083), .A2(n1081), .ZN(n1080) );
  MUX2ND0 U1229 ( .I0(N59), .I1(mantissa_ab[14]), .S(n553), .ZN(n1121) );
  MUX2D0 U1230 ( .I0(mantissa_ab[13]), .I1(n747), .S(n593), .Z(
        comp_mantissa_ab[13]) );
  XNR2D0 U1231 ( .A1(n1134), .A2(n1122), .ZN(n747) );
  MUX2ND0 U1232 ( .I0(mantissa_ab[13]), .I1(N58), .S(n904), .ZN(n1122) );
  NR2D0 U1233 ( .A1(n1113), .A2(n549), .ZN(n1134) );
  AN2D0 U1234 ( .A1(n1135), .A2(n1117), .Z(n1113) );
  AN3D0 U1235 ( .A1(n1111), .A2(n1136), .A3(n1137), .Z(n1117) );
  MUX2D0 U1236 ( .I0(mantissa_ab[12]), .I1(n758), .S(n593), .Z(
        comp_mantissa_ab[12]) );
  XNR2D0 U1237 ( .A1(n1138), .A2(n1111), .ZN(n758) );
  MUX2ND0 U1238 ( .I0(mantissa_ab[12]), .I1(N57), .S(n904), .ZN(n1111) );
  NR2D0 U1239 ( .A1(n1109), .A2(n549), .ZN(n1138) );
  CKND0 U1240 ( .I(sign_ab), .ZN(n549) );
  MUX2D0 U1241 ( .I0(mantissa_ab[11]), .I1(n771), .S(n593), .Z(
        comp_mantissa_ab[11]) );
  INR2D0 U1242 ( .A1(n1139), .B1(n1109), .ZN(n771) );
  INR2D0 U1243 ( .A1(n1137), .B1(n1140), .ZN(n1109) );
  MUX2ND0 U1244 ( .I0(n1137), .I1(n1141), .S(sign_ab), .ZN(n1139) );
  INR2D0 U1245 ( .A1(n1140), .B1(n1137), .ZN(n1141) );
  MUX2ND0 U1246 ( .I0(N56), .I1(mantissa_ab[11]), .S(n553), .ZN(n1137) );
  MUX2D0 U1247 ( .I0(mantissa_ab[10]), .I1(n782), .S(n593), .Z(
        comp_mantissa_ab[10]) );
  CKND0 U1248 ( .I(n823), .ZN(n782) );
  CKND2D0 U1249 ( .A1(n1142), .A2(n1140), .ZN(n823) );
  CKND2D0 U1250 ( .A1(n1135), .A2(n1136), .ZN(n1140) );
  MUX2ND0 U1251 ( .I0(n1136), .I1(n1143), .S(sign_ab), .ZN(n1142) );
  NR2D0 U1252 ( .A1(n1135), .A2(n1136), .ZN(n1143) );
  AN3D0 U1253 ( .A1(n1083), .A2(n1064), .A3(n1123), .Z(n1135) );
  AN4D0 U1254 ( .A1(n1067), .A2(n1071), .A3(n1076), .A4(n1081), .Z(n1123) );
  MUX2ND0 U1255 ( .I0(N50), .I1(mantissa_ab[5]), .S(n553), .ZN(n1081) );
  MUX2ND0 U1256 ( .I0(N51), .I1(mantissa_ab[6]), .S(n553), .ZN(n1076) );
  MUX2ND0 U1257 ( .I0(N52), .I1(mantissa_ab[7]), .S(n553), .ZN(n1071) );
  MUX2ND0 U1258 ( .I0(mantissa_ab[8]), .I1(N53), .S(n904), .ZN(n1067) );
  MUX2ND0 U1259 ( .I0(mantissa_ab[9]), .I1(N54), .S(n904), .ZN(n1064) );
  CKND0 U1260 ( .I(n1085), .ZN(n1083) );
  CKND2D0 U1261 ( .A1(n1088), .A2(n1086), .ZN(n1085) );
  MUX2ND0 U1262 ( .I0(N49), .I1(mantissa_ab[4]), .S(n553), .ZN(n1086) );
  CKND0 U1263 ( .I(n1090), .ZN(n1088) );
  CKND2D0 U1264 ( .A1(n1093), .A2(n1091), .ZN(n1090) );
  MUX2ND0 U1265 ( .I0(N48), .I1(mantissa_ab[3]), .S(n553), .ZN(n1091) );
  INR2D0 U1266 ( .A1(n1095), .B1(n1097), .ZN(n1093) );
  CKND2D0 U1267 ( .A1(n1106), .A2(n844), .ZN(n1097) );
  MUX2ND0 U1268 ( .I0(mantissa_ab[1]), .I1(N46), .S(n904), .ZN(n1106) );
  MUX2ND0 U1269 ( .I0(mantissa_ab[2]), .I1(N47), .S(n904), .ZN(n1095) );
  MUX2ND0 U1270 ( .I0(N55), .I1(mantissa_ab[10]), .S(n553), .ZN(n1136) );
  MUX2ND0 U1271 ( .I0(n844), .I1(n1144), .S(fma_byp), .ZN(comp_mantissa_ab[0])
         );
  CKND0 U1272 ( .I(mantissa_ab[0]), .ZN(n1144) );
  MUX2ND0 U1273 ( .I0(mantissa_ab[0]), .I1(N45), .S(n904), .ZN(n844) );
  CKND0 U1274 ( .I(n553), .ZN(n904) );
  CKND2D0 U1275 ( .A1(exp_ab_less), .A2(n547), .ZN(n553) );
  CKND0 U1276 ( .I(exp_ab_greater), .ZN(n547) );
  ND4D0 U1277 ( .A1(n903), .A2(n901), .A3(n1145), .A4(n899), .ZN(N800) );
  CKND0 U1278 ( .I(exp_ab[2]), .ZN(n899) );
  NR2D0 U1279 ( .A1(exp_ab[4]), .A2(exp_ab[3]), .ZN(n1145) );
  CKND0 U1280 ( .I(exp_ab[1]), .ZN(n901) );
  CKND0 U1281 ( .I(exp_ab[0]), .ZN(n903) );
endmodule

