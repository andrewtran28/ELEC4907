
module arbiter ( clk, rst, fifo_empty, fifo_0_snoop, fifo_1_snoop, 
        fifo_2_snoop, fifo_3_snoop, fifo_4_snoop, fifo_5_snoop, fifo_6_snoop, 
        fifo_7_snoop, router_ready, ready, fifo_rd, fifo_0_ptr, fifo_1_ptr, 
        fifo_2_ptr, fifo_3_ptr, fifo_4_ptr, fifo_5_ptr, fifo_6_ptr, fifo_7_ptr
 );
  input [7:0] fifo_empty;
  input [31:0] fifo_0_snoop;
  input [31:0] fifo_1_snoop;
  input [31:0] fifo_2_snoop;
  input [31:0] fifo_3_snoop;
  input [31:0] fifo_4_snoop;
  input [31:0] fifo_5_snoop;
  input [31:0] fifo_6_snoop;
  input [31:0] fifo_7_snoop;
  output [2:0] fifo_0_ptr;
  output [2:0] fifo_1_ptr;
  output [2:0] fifo_2_ptr;
  output [2:0] fifo_3_ptr;
  output [2:0] fifo_4_ptr;
  output [2:0] fifo_5_ptr;
  output [2:0] fifo_6_ptr;
  output [2:0] fifo_7_ptr;
  input clk, rst, router_ready;
  output ready, fifo_rd;
  wire   N3079, N3080, N3081, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616;

  DFQD1 \fifo_7_ptr_reg[2]  ( .D(n2895), .CP(clk), .Q(fifo_7_ptr[2]) );
  DFQD1 \fifo_7_ptr_reg[1]  ( .D(n2894), .CP(clk), .Q(fifo_7_ptr[1]) );
  DFQD1 \fifo_7_ptr_reg[0]  ( .D(n2893), .CP(clk), .Q(fifo_7_ptr[0]) );
  DFQD1 \fifo_2_ptr_reg[2]  ( .D(n2892), .CP(clk), .Q(fifo_2_ptr[2]) );
  DFQD1 \fifo_2_ptr_reg[1]  ( .D(n2891), .CP(clk), .Q(fifo_2_ptr[1]) );
  DFQD1 \fifo_2_ptr_reg[0]  ( .D(n2890), .CP(clk), .Q(fifo_2_ptr[0]) );
  DFQD1 \fifo_1_ptr_reg[2]  ( .D(n2889), .CP(clk), .Q(fifo_1_ptr[2]) );
  DFQD1 \fifo_1_ptr_reg[1]  ( .D(n2888), .CP(clk), .Q(fifo_1_ptr[1]) );
  DFQD1 \fifo_1_ptr_reg[0]  ( .D(n2887), .CP(clk), .Q(fifo_1_ptr[0]) );
  EDFQD1 \fifo_0_ptr_reg[2]  ( .D(N3081), .E(n2896), .CP(clk), .Q(
        fifo_0_ptr[2]) );
  EDFQD1 \fifo_0_ptr_reg[1]  ( .D(N3080), .E(n2896), .CP(clk), .Q(
        fifo_0_ptr[1]) );
  EDFQD1 \fifo_0_ptr_reg[0]  ( .D(N3079), .E(n2896), .CP(clk), .Q(
        fifo_0_ptr[0]) );
  DFQD1 \fifo_3_ptr_reg[2]  ( .D(n2886), .CP(clk), .Q(fifo_3_ptr[2]) );
  DFQD1 \fifo_3_ptr_reg[1]  ( .D(n2885), .CP(clk), .Q(fifo_3_ptr[1]) );
  DFQD1 \fifo_3_ptr_reg[0]  ( .D(n2884), .CP(clk), .Q(fifo_3_ptr[0]) );
  DFQD1 \fifo_5_ptr_reg[2]  ( .D(n2883), .CP(clk), .Q(fifo_5_ptr[2]) );
  DFQD1 \fifo_5_ptr_reg[1]  ( .D(n2882), .CP(clk), .Q(fifo_5_ptr[1]) );
  DFQD1 \fifo_5_ptr_reg[0]  ( .D(n2881), .CP(clk), .Q(fifo_5_ptr[0]) );
  DFQD1 \fifo_4_ptr_reg[2]  ( .D(n2880), .CP(clk), .Q(fifo_4_ptr[2]) );
  DFQD1 \fifo_4_ptr_reg[1]  ( .D(n2879), .CP(clk), .Q(fifo_4_ptr[1]) );
  DFQD1 \fifo_4_ptr_reg[0]  ( .D(n2878), .CP(clk), .Q(fifo_4_ptr[0]) );
  DFQD1 \fifo_6_ptr_reg[2]  ( .D(n2877), .CP(clk), .Q(fifo_6_ptr[2]) );
  DFQD1 \fifo_6_ptr_reg[1]  ( .D(n2876), .CP(clk), .Q(fifo_6_ptr[1]) );
  DFQD1 \fifo_6_ptr_reg[0]  ( .D(n2875), .CP(clk), .Q(fifo_6_ptr[0]) );
  TIEH U2903 ( .Z(ready) );
  MUX2D0 U2904 ( .I0(fifo_7_ptr[2]), .I1(n2897), .S(n2898), .Z(n2895) );
  CKND2D0 U2905 ( .A1(n2899), .A2(n2900), .ZN(n2897) );
  AOI221D0 U2906 ( .A1(n2901), .A2(n2902), .B1(n2903), .B2(n2904), .C(n2905), 
        .ZN(n2900) );
  OAI22D0 U2907 ( .A1(n2906), .A2(n2907), .B1(n2908), .B2(n2909), .ZN(n2905)
         );
  AOI222D0 U2908 ( .A1(n2910), .A2(n2911), .B1(n2912), .B2(n2913), .C1(n2914), 
        .C2(n2915), .ZN(n2899) );
  MUX2D0 U2909 ( .I0(fifo_7_ptr[1]), .I1(n2916), .S(n2898), .Z(n2894) );
  CKND2D0 U2910 ( .A1(n2917), .A2(n2918), .ZN(n2916) );
  AOI221D0 U2911 ( .A1(n2901), .A2(n2919), .B1(n2903), .B2(n2920), .C(n2921), 
        .ZN(n2918) );
  OAI22D0 U2912 ( .A1(n2922), .A2(n2907), .B1(n2923), .B2(n2909), .ZN(n2921)
         );
  AOI222D0 U2913 ( .A1(n2910), .A2(n2924), .B1(n2912), .B2(n2925), .C1(n2914), 
        .C2(n2926), .ZN(n2917) );
  MUX2D0 U2914 ( .I0(fifo_7_ptr[0]), .I1(n2927), .S(n2898), .Z(n2893) );
  OA31D0 U2915 ( .A1(n2928), .A2(n2912), .A3(n2929), .B(n2896), .Z(n2898) );
  OAI31D0 U2916 ( .A1(n2930), .A2(n2931), .A3(n2932), .B(n2933), .ZN(n2929) );
  ND4D0 U2917 ( .A1(n2934), .A2(n2909), .A3(n2907), .A4(n2935), .ZN(n2928) );
  CKND2D0 U2918 ( .A1(n2936), .A2(n2937), .ZN(n2927) );
  AOI221D0 U2919 ( .A1(n2901), .A2(n2938), .B1(n2903), .B2(n2939), .C(n2940), 
        .ZN(n2937) );
  OAI22D0 U2920 ( .A1(n2941), .A2(n2907), .B1(n2942), .B2(n2909), .ZN(n2940)
         );
  ND4D0 U2921 ( .A1(n2943), .A2(n2944), .A3(n2945), .A4(n2946), .ZN(n2909) );
  CKND2D0 U2922 ( .A1(n2947), .A2(n2944), .ZN(n2907) );
  CKND0 U2923 ( .I(n2934), .ZN(n2903) );
  CKND2D0 U2924 ( .A1(n2948), .A2(n2949), .ZN(n2934) );
  CKND0 U2925 ( .I(n2932), .ZN(n2901) );
  OAI31D0 U2926 ( .A1(n2950), .A2(n2951), .A3(n2952), .B(n2949), .ZN(n2932) );
  OA31D0 U2927 ( .A1(n2953), .A2(n2954), .A3(n2955), .B(n2956), .Z(n2949) );
  AOI222D0 U2928 ( .A1(n2910), .A2(n2957), .B1(n2912), .B2(n2958), .C1(n2914), 
        .C2(n2959), .ZN(n2936) );
  CKND0 U2929 ( .I(n2933), .ZN(n2914) );
  CKND2D0 U2930 ( .A1(n2960), .A2(n2961), .ZN(n2933) );
  AN2D0 U2931 ( .A1(n2962), .A2(n2956), .Z(n2912) );
  OA211D0 U2932 ( .A1(n2963), .A2(n2964), .B(n2946), .C(n2944), .Z(n2956) );
  OA31D0 U2933 ( .A1(n2965), .A2(n2966), .A3(n2967), .B(n2961), .Z(n2944) );
  ND3D0 U2934 ( .A1(n2968), .A2(n2969), .A3(n2970), .ZN(n2961) );
  ND3D0 U2935 ( .A1(n2971), .A2(n2972), .A3(n2973), .ZN(n2946) );
  NR2D0 U2936 ( .A1(n2974), .A2(n2945), .ZN(n2963) );
  MUX2D0 U2937 ( .I0(fifo_2_ptr[2]), .I1(n2975), .S(n2976), .Z(n2892) );
  CKND2D0 U2938 ( .A1(n2977), .A2(n2978), .ZN(n2975) );
  AOI221D0 U2939 ( .A1(n2979), .A2(n2902), .B1(n2980), .B2(n2904), .C(n2981), 
        .ZN(n2978) );
  OAI22D0 U2940 ( .A1(n2906), .A2(n2982), .B1(n2908), .B2(n2983), .ZN(n2981)
         );
  AOI222D0 U2941 ( .A1(n2984), .A2(n2911), .B1(n2985), .B2(n2913), .C1(n2986), 
        .C2(n2915), .ZN(n2977) );
  MUX2D0 U2942 ( .I0(fifo_2_ptr[1]), .I1(n2987), .S(n2976), .Z(n2891) );
  CKND2D0 U2943 ( .A1(n2988), .A2(n2989), .ZN(n2987) );
  AOI221D0 U2944 ( .A1(n2979), .A2(n2919), .B1(n2980), .B2(n2920), .C(n2990), 
        .ZN(n2989) );
  OAI22D0 U2945 ( .A1(n2922), .A2(n2982), .B1(n2923), .B2(n2983), .ZN(n2990)
         );
  AOI222D0 U2946 ( .A1(n2984), .A2(n2924), .B1(n2985), .B2(n2925), .C1(n2986), 
        .C2(n2926), .ZN(n2988) );
  MUX2D0 U2947 ( .I0(fifo_2_ptr[0]), .I1(n2991), .S(n2976), .Z(n2890) );
  OA31D0 U2948 ( .A1(n2992), .A2(n2986), .A3(n2993), .B(n2896), .Z(n2976) );
  CKND2D0 U2949 ( .A1(n2994), .A2(n2995), .ZN(n2993) );
  OAI211D0 U2950 ( .A1(n2996), .A2(n2997), .B(n2998), .C(n2999), .ZN(n2992) );
  ND4D0 U2951 ( .A1(n2979), .A2(n3000), .A3(n2931), .A4(n3001), .ZN(n2998) );
  NR2D0 U2952 ( .A1(n3002), .A2(n3003), .ZN(n2996) );
  CKND2D0 U2953 ( .A1(n3004), .A2(n3005), .ZN(n2991) );
  AOI221D0 U2954 ( .A1(n2979), .A2(n2938), .B1(n2980), .B2(n2939), .C(n3006), 
        .ZN(n3005) );
  OAI22D0 U2955 ( .A1(n2941), .A2(n2982), .B1(n2942), .B2(n2983), .ZN(n3006)
         );
  CKND2D0 U2956 ( .A1(n3003), .A2(n3007), .ZN(n2983) );
  AN2D0 U2957 ( .A1(n3008), .A2(n3009), .Z(n3003) );
  CKND2D0 U2958 ( .A1(n3002), .A2(n3007), .ZN(n2982) );
  CKND0 U2959 ( .I(n2994), .ZN(n2980) );
  CKND2D0 U2960 ( .A1(n3010), .A2(n3011), .ZN(n2994) );
  OA21D0 U2961 ( .A1(n3012), .A2(n3013), .B(n3011), .Z(n2979) );
  OA31D0 U2962 ( .A1(n3014), .A2(n3015), .A3(n3016), .B(n3017), .Z(n3011) );
  AOI222D0 U2963 ( .A1(n2984), .A2(n2957), .B1(n2985), .B2(n2958), .C1(n2986), 
        .C2(n2959), .ZN(n3004) );
  AN2D0 U2964 ( .A1(n3018), .A2(n3019), .Z(n2986) );
  CKND0 U2965 ( .I(n2999), .ZN(n2985) );
  CKND2D0 U2966 ( .A1(n3020), .A2(n3017), .ZN(n2999) );
  OA211D0 U2967 ( .A1(n3021), .A2(n3022), .B(n3009), .C(n3007), .Z(n3017) );
  CKND0 U2968 ( .I(n2997), .ZN(n3007) );
  OAI31D0 U2969 ( .A1(n3023), .A2(n3024), .A3(n3025), .B(n3018), .ZN(n2997) );
  CKND2D0 U2970 ( .A1(n3026), .A2(n3027), .ZN(n3018) );
  CKND2D0 U2971 ( .A1(n3028), .A2(n3029), .ZN(n3009) );
  MUX2D0 U2972 ( .I0(fifo_1_ptr[2]), .I1(n3030), .S(n3031), .Z(n2889) );
  CKND2D0 U2973 ( .A1(n3032), .A2(n3033), .ZN(n3030) );
  AOI221D0 U2974 ( .A1(n3034), .A2(n2902), .B1(n3035), .B2(n2904), .C(n3036), 
        .ZN(n3033) );
  OAI22D0 U2975 ( .A1(n2906), .A2(n3037), .B1(n2908), .B2(n3038), .ZN(n3036)
         );
  AOI222D0 U2976 ( .A1(n3039), .A2(n2911), .B1(n3040), .B2(n2913), .C1(n3041), 
        .C2(n2915), .ZN(n3032) );
  MUX2D0 U2977 ( .I0(fifo_1_ptr[1]), .I1(n3042), .S(n3031), .Z(n2888) );
  CKND2D0 U2978 ( .A1(n3043), .A2(n3044), .ZN(n3042) );
  AOI221D0 U2979 ( .A1(n3034), .A2(n2919), .B1(n3035), .B2(n2920), .C(n3045), 
        .ZN(n3044) );
  OAI22D0 U2980 ( .A1(n2922), .A2(n3037), .B1(n2923), .B2(n3038), .ZN(n3045)
         );
  AOI222D0 U2981 ( .A1(n3039), .A2(n2924), .B1(n3040), .B2(n2925), .C1(n3041), 
        .C2(n2926), .ZN(n3043) );
  MUX2D0 U2982 ( .I0(fifo_1_ptr[0]), .I1(n3046), .S(n3031), .Z(n2887) );
  OA31D0 U2983 ( .A1(n3047), .A2(n3041), .A3(n3048), .B(n2896), .Z(n3031) );
  CKND2D0 U2984 ( .A1(n3049), .A2(n3027), .ZN(n3048) );
  OAI211D0 U2985 ( .A1(n3050), .A2(n3051), .B(n3052), .C(n3053), .ZN(n3047) );
  ND4D0 U2986 ( .A1(n3054), .A2(n3034), .A3(n3000), .A4(n3055), .ZN(n3052) );
  NR2D0 U2987 ( .A1(n3056), .A2(n3057), .ZN(n3050) );
  CKND2D0 U2988 ( .A1(n3058), .A2(n3059), .ZN(n3046) );
  AOI221D0 U2989 ( .A1(n3034), .A2(n2938), .B1(n3035), .B2(n2939), .C(n3060), 
        .ZN(n3059) );
  OAI22D0 U2990 ( .A1(n2941), .A2(n3037), .B1(n2942), .B2(n3038), .ZN(n3060)
         );
  CKND2D0 U2991 ( .A1(n3057), .A2(n3061), .ZN(n3038) );
  AN2D0 U2992 ( .A1(n3021), .A2(n3062), .Z(n3057) );
  CKND2D0 U2993 ( .A1(n3056), .A2(n3061), .ZN(n3037) );
  CKND0 U2994 ( .I(n3049), .ZN(n3035) );
  CKND2D0 U2995 ( .A1(n3012), .A2(n3063), .ZN(n3049) );
  OA21D0 U2996 ( .A1(n3010), .A2(n3013), .B(n3063), .Z(n3034) );
  OA31D0 U2997 ( .A1(n3014), .A2(n3020), .A3(n3016), .B(n3064), .Z(n3063) );
  OR4D0 U2998 ( .A1(n2955), .A2(n2962), .A3(n2954), .A4(n3065), .Z(n3014) );
  ND4D0 U2999 ( .A1(n3066), .A2(n3067), .A3(n3068), .A4(n3069), .ZN(n3013) );
  NR3D0 U3000 ( .A1(n2952), .A2(n2951), .A3(n2948), .ZN(n3069) );
  AOI222D0 U3001 ( .A1(n3039), .A2(n2957), .B1(n3040), .B2(n2958), .C1(n3041), 
        .C2(n2959), .ZN(n3058) );
  AN2D0 U3002 ( .A1(n3024), .A2(n3070), .Z(n3041) );
  CKND0 U3003 ( .I(n3053), .ZN(n3040) );
  CKND2D0 U3004 ( .A1(n3015), .A2(n3064), .ZN(n3053) );
  OA211D0 U3005 ( .A1(n3008), .A2(n3022), .B(n3062), .C(n3061), .Z(n3064) );
  CKND0 U3006 ( .I(n3051), .ZN(n3061) );
  OAI31D0 U3007 ( .A1(n3023), .A2(n3019), .A3(n3025), .B(n3070), .ZN(n3051) );
  CKND2D0 U3008 ( .A1(n3026), .A2(n2995), .ZN(n3070) );
  INR4D0 U3009 ( .A1(n3071), .B1(n2910), .B2(n3072), .B3(n3073), .ZN(n3026) );
  NR3D0 U3010 ( .A1(n3074), .A2(n3075), .A3(n3076), .ZN(n3071) );
  OR4D0 U3011 ( .A1(n2967), .A2(n2960), .A3(n2966), .A4(n3077), .Z(n3023) );
  CKND2D0 U3012 ( .A1(n3028), .A2(n3078), .ZN(n3062) );
  INR4D0 U3013 ( .A1(n3079), .B1(n2947), .B2(n3080), .B3(n3081), .ZN(n3028) );
  NR3D0 U3014 ( .A1(n3082), .A2(n3083), .A3(n3084), .ZN(n3079) );
  ND4D0 U3015 ( .A1(n3085), .A2(n3086), .A3(n3087), .A4(n2974), .ZN(n3022) );
  MUX2D0 U3016 ( .I0(fifo_3_ptr[2]), .I1(n3088), .S(n3089), .Z(n2886) );
  CKND2D0 U3017 ( .A1(n3090), .A2(n3091), .ZN(n3088) );
  AOI221D0 U3018 ( .A1(n3092), .A2(n2902), .B1(n3093), .B2(n2904), .C(n3094), 
        .ZN(n3091) );
  OAI22D0 U3019 ( .A1(n2906), .A2(n3095), .B1(n2908), .B2(n3096), .ZN(n3094)
         );
  AOI222D0 U3020 ( .A1(n3075), .A2(n2911), .B1(n3097), .B2(n2913), .C1(n3098), 
        .C2(n2915), .ZN(n3090) );
  MUX2D0 U3021 ( .I0(fifo_3_ptr[1]), .I1(n3099), .S(n3089), .Z(n2885) );
  CKND2D0 U3022 ( .A1(n3100), .A2(n3101), .ZN(n3099) );
  AOI221D0 U3023 ( .A1(n3092), .A2(n2919), .B1(n3093), .B2(n2920), .C(n3102), 
        .ZN(n3101) );
  OAI22D0 U3024 ( .A1(n2922), .A2(n3095), .B1(n2923), .B2(n3096), .ZN(n3102)
         );
  AOI222D0 U3025 ( .A1(n3075), .A2(n2924), .B1(n3097), .B2(n2925), .C1(n3098), 
        .C2(n2926), .ZN(n3100) );
  MUX2D0 U3026 ( .I0(fifo_3_ptr[0]), .I1(n3103), .S(n3089), .Z(n2884) );
  OA31D0 U3027 ( .A1(n3104), .A2(n3097), .A3(n3105), .B(n2896), .Z(n3089) );
  OAI31D0 U3028 ( .A1(n3106), .A2(n3107), .A3(n3108), .B(n3109), .ZN(n3105) );
  CKND2D0 U3029 ( .A1(n3055), .A2(n3001), .ZN(n3106) );
  ND4D0 U3030 ( .A1(n3110), .A2(n3096), .A3(n3095), .A4(n3111), .ZN(n3104) );
  CKND2D0 U3031 ( .A1(n3112), .A2(n3113), .ZN(n3103) );
  AOI221D0 U3032 ( .A1(n3092), .A2(n2938), .B1(n3093), .B2(n2939), .C(n3114), 
        .ZN(n3113) );
  OAI22D0 U3033 ( .A1(n2941), .A2(n3095), .B1(n2942), .B2(n3096), .ZN(n3114)
         );
  ND3D0 U3034 ( .A1(n3115), .A2(n3116), .A3(n3117), .ZN(n3096) );
  CKND2D0 U3035 ( .A1(n3083), .A2(n3115), .ZN(n3095) );
  CKND0 U3036 ( .I(n3110), .ZN(n3093) );
  CKND2D0 U3037 ( .A1(n3118), .A2(n3119), .ZN(n3110) );
  CKND0 U3038 ( .I(n3108), .ZN(n3092) );
  OAI31D0 U3039 ( .A1(n3120), .A2(n3121), .A3(n3122), .B(n3119), .ZN(n3108) );
  OA31D0 U3040 ( .A1(n3123), .A2(n3065), .A3(n3124), .B(n3125), .Z(n3119) );
  AOI222D0 U3041 ( .A1(n3075), .A2(n2957), .B1(n3097), .B2(n2958), .C1(n3098), 
        .C2(n2959), .ZN(n3112) );
  CKND0 U3042 ( .I(n3109), .ZN(n3098) );
  CKND2D0 U3043 ( .A1(n3126), .A2(n3127), .ZN(n3109) );
  AN2D0 U3044 ( .A1(n3128), .A2(n3125), .Z(n3097) );
  OA211D0 U3045 ( .A1(n3129), .A2(n3130), .B(n3116), .C(n3115), .Z(n3125) );
  OA31D0 U3046 ( .A1(n3131), .A2(n3077), .A3(n3132), .B(n3127), .Z(n3115) );
  ND3D0 U3047 ( .A1(n3133), .A2(n3134), .A3(n3135), .ZN(n3127) );
  ND3D0 U3048 ( .A1(n3136), .A2(n3137), .A3(n3138), .ZN(n3116) );
  MUX2D0 U3049 ( .I0(fifo_5_ptr[2]), .I1(n3139), .S(n3140), .Z(n2883) );
  CKND2D0 U3050 ( .A1(n3141), .A2(n3142), .ZN(n3139) );
  AOI221D0 U3051 ( .A1(n3143), .A2(n2902), .B1(n3144), .B2(n2904), .C(n3145), 
        .ZN(n3142) );
  OAI22D0 U3052 ( .A1(n2906), .A2(n3146), .B1(n2908), .B2(n3147), .ZN(n3145)
         );
  AOI222D0 U3053 ( .A1(n3073), .A2(n2911), .B1(n3148), .B2(n2913), .C1(n3149), 
        .C2(n2915), .ZN(n3141) );
  MUX2D0 U3054 ( .I0(fifo_5_ptr[1]), .I1(n3150), .S(n3140), .Z(n2882) );
  CKND2D0 U3055 ( .A1(n3151), .A2(n3152), .ZN(n3150) );
  AOI221D0 U3056 ( .A1(n3143), .A2(n2919), .B1(n3144), .B2(n2920), .C(n3153), 
        .ZN(n3152) );
  OAI22D0 U3057 ( .A1(n2922), .A2(n3146), .B1(n2923), .B2(n3147), .ZN(n3153)
         );
  AOI222D0 U3058 ( .A1(n3073), .A2(n2924), .B1(n3148), .B2(n2925), .C1(n3149), 
        .C2(n2926), .ZN(n3151) );
  MUX2D0 U3059 ( .I0(fifo_5_ptr[0]), .I1(n3154), .S(n3140), .Z(n2881) );
  AN2D0 U3060 ( .A1(n2896), .A2(n3155), .Z(n3140) );
  ND4D0 U3061 ( .A1(n3156), .A2(n2968), .A3(n3157), .A4(n3158), .ZN(n3155) );
  AOI211D0 U3062 ( .A1(n3159), .A2(n3160), .B(n3148), .C(n3161), .ZN(n3158) );
  NR4D0 U3063 ( .A1(n3000), .A2(n2931), .A3(n3001), .A4(n3162), .ZN(n3161) );
  CKND2D0 U3064 ( .A1(n3163), .A2(n2971), .ZN(n3160) );
  CKND2D0 U3065 ( .A1(n3164), .A2(n3165), .ZN(n3154) );
  AOI221D0 U3066 ( .A1(n3143), .A2(n2938), .B1(n3144), .B2(n2939), .C(n3166), 
        .ZN(n3165) );
  OAI22D0 U3067 ( .A1(n2941), .A2(n3146), .B1(n2942), .B2(n3147), .ZN(n3166)
         );
  IND2D0 U3068 ( .A1(n3163), .B1(n3159), .ZN(n3147) );
  CKND2D0 U3069 ( .A1(n3167), .A2(n3168), .ZN(n3163) );
  CKND2D0 U3070 ( .A1(n3081), .A2(n3159), .ZN(n3146) );
  CKND0 U3071 ( .I(n3156), .ZN(n3144) );
  CKND2D0 U3072 ( .A1(n2952), .A2(n3169), .ZN(n3156) );
  CKND0 U3073 ( .I(n3162), .ZN(n3143) );
  OAI31D0 U3074 ( .A1(n2950), .A2(n2951), .A3(n2948), .B(n3169), .ZN(n3162) );
  OA31D0 U3075 ( .A1(n2953), .A2(n2954), .A3(n2962), .B(n3170), .Z(n3169) );
  AOI222D0 U3076 ( .A1(n3073), .A2(n2957), .B1(n3148), .B2(n2958), .C1(n3149), 
        .C2(n2959), .ZN(n3164) );
  CKND0 U3077 ( .I(n3157), .ZN(n3149) );
  CKND2D0 U3078 ( .A1(n2967), .A2(n3171), .ZN(n3157) );
  AN2D0 U3079 ( .A1(n2955), .A2(n3170), .Z(n3148) );
  OA211D0 U3080 ( .A1(n2943), .A2(n3172), .B(n3168), .C(n3159), .Z(n3170) );
  OA31D0 U3081 ( .A1(n2965), .A2(n2966), .A3(n2960), .B(n3171), .Z(n3159) );
  ND3D0 U3082 ( .A1(n2935), .A2(n2969), .A3(n2970), .ZN(n3171) );
  ND3D0 U3083 ( .A1(n3173), .A2(n2972), .A3(n2973), .ZN(n3168) );
  CKND0 U3084 ( .I(n3174), .ZN(n3172) );
  MUX2D0 U3085 ( .I0(fifo_4_ptr[2]), .I1(n3175), .S(n3176), .Z(n2880) );
  CKND2D0 U3086 ( .A1(n3177), .A2(n3178), .ZN(n3175) );
  AOI221D0 U3087 ( .A1(n3179), .A2(n2902), .B1(n3180), .B2(n2904), .C(n3181), 
        .ZN(n3178) );
  OAI22D0 U3088 ( .A1(n2906), .A2(n3182), .B1(n2908), .B2(n3183), .ZN(n3181)
         );
  AOI222D0 U3089 ( .A1(n3076), .A2(n2911), .B1(n3184), .B2(n2913), .C1(n3185), 
        .C2(n2915), .ZN(n3177) );
  MUX2D0 U3090 ( .I0(fifo_4_ptr[1]), .I1(n3186), .S(n3176), .Z(n2879) );
  CKND2D0 U3091 ( .A1(n3187), .A2(n3188), .ZN(n3186) );
  AOI221D0 U3092 ( .A1(n3179), .A2(n2919), .B1(n3180), .B2(n2920), .C(n3189), 
        .ZN(n3188) );
  OAI22D0 U3093 ( .A1(n2922), .A2(n3182), .B1(n2923), .B2(n3183), .ZN(n3189)
         );
  AOI222D0 U3094 ( .A1(n3076), .A2(n2924), .B1(n3184), .B2(n2925), .C1(n3185), 
        .C2(n2926), .ZN(n3187) );
  MUX2D0 U3095 ( .I0(fifo_4_ptr[0]), .I1(n3190), .S(n3176), .Z(n2878) );
  OA31D0 U3096 ( .A1(n3191), .A2(n3184), .A3(n3192), .B(n2896), .Z(n3176) );
  OAI31D0 U3097 ( .A1(n3193), .A2(n3001), .A3(n3194), .B(n3195), .ZN(n3192) );
  CKND2D0 U3098 ( .A1(n2931), .A2(n3107), .ZN(n3193) );
  CKND0 U3099 ( .I(n3055), .ZN(n2931) );
  ND4D0 U3100 ( .A1(n3196), .A2(n3183), .A3(n3182), .A4(n3134), .ZN(n3191) );
  CKND2D0 U3101 ( .A1(n3197), .A2(n3198), .ZN(n3190) );
  AOI221D0 U3102 ( .A1(n3179), .A2(n2938), .B1(n3180), .B2(n2939), .C(n3199), 
        .ZN(n3198) );
  OAI22D0 U3103 ( .A1(n2941), .A2(n3182), .B1(n2942), .B2(n3183), .ZN(n3199)
         );
  ND3D0 U3104 ( .A1(n3200), .A2(n3201), .A3(n3129), .ZN(n3183) );
  CKND2D0 U3105 ( .A1(n3084), .A2(n3200), .ZN(n3182) );
  CKND0 U3106 ( .I(n3196), .ZN(n3180) );
  CKND2D0 U3107 ( .A1(n3121), .A2(n3202), .ZN(n3196) );
  CKND0 U3108 ( .I(n3066), .ZN(n3121) );
  CKND0 U3109 ( .I(n3194), .ZN(n3179) );
  OAI31D0 U3110 ( .A1(n3120), .A2(n3118), .A3(n3122), .B(n3202), .ZN(n3194) );
  OA31D0 U3111 ( .A1(n3123), .A2(n3065), .A3(n3128), .B(n3203), .Z(n3202) );
  CKND0 U3112 ( .I(n3068), .ZN(n3122) );
  CKND0 U3113 ( .I(n3067), .ZN(n3118) );
  CKND0 U3114 ( .I(n3204), .ZN(n3120) );
  AOI222D0 U3115 ( .A1(n3076), .A2(n2957), .B1(n3184), .B2(n2958), .C1(n3185), 
        .C2(n2959), .ZN(n3197) );
  CKND0 U3116 ( .I(n3195), .ZN(n3185) );
  CKND2D0 U3117 ( .A1(n3132), .A2(n3205), .ZN(n3195) );
  AN2D0 U3118 ( .A1(n3124), .A2(n3203), .Z(n3184) );
  OA211D0 U3119 ( .A1(n3117), .A2(n3130), .B(n3201), .C(n3200), .Z(n3203) );
  OA31D0 U3120 ( .A1(n3131), .A2(n3077), .A3(n3126), .B(n3205), .Z(n3200) );
  ND3D0 U3121 ( .A1(n3133), .A2(n3111), .A3(n3135), .ZN(n3205) );
  ND3D0 U3122 ( .A1(n3136), .A2(n3206), .A3(n3138), .ZN(n3201) );
  CKND2D0 U3123 ( .A1(n3207), .A2(n3087), .ZN(n3130) );
  MUX2D0 U3124 ( .I0(fifo_6_ptr[2]), .I1(n3208), .S(n3209), .Z(n2877) );
  CKND2D0 U3125 ( .A1(n3210), .A2(n3211), .ZN(n3208) );
  AOI221D0 U3126 ( .A1(n3212), .A2(n2902), .B1(n3213), .B2(n2904), .C(n3214), 
        .ZN(n3211) );
  OAI22D0 U3127 ( .A1(n2906), .A2(n3215), .B1(n2908), .B2(n3216), .ZN(n3214)
         );
  CKND0 U3128 ( .I(n3217), .ZN(n2908) );
  AOI222D0 U3129 ( .A1(n3072), .A2(n2911), .B1(n3218), .B2(n2913), .C1(n3219), 
        .C2(n2915), .ZN(n3210) );
  MUX2D0 U3130 ( .I0(fifo_6_ptr[1]), .I1(n3220), .S(n3209), .Z(n2876) );
  CKND2D0 U3131 ( .A1(n3221), .A2(n3222), .ZN(n3220) );
  AOI221D0 U3132 ( .A1(n3212), .A2(n2919), .B1(n3213), .B2(n2920), .C(n3223), 
        .ZN(n3222) );
  OAI22D0 U3133 ( .A1(n2922), .A2(n3215), .B1(n2923), .B2(n3216), .ZN(n3223)
         );
  CKND0 U3134 ( .I(n3224), .ZN(n2923) );
  AOI222D0 U3135 ( .A1(n3072), .A2(n2924), .B1(n3218), .B2(n2925), .C1(n3219), 
        .C2(n2926), .ZN(n3221) );
  MUX2D0 U3136 ( .I0(fifo_6_ptr[0]), .I1(n3225), .S(n3209), .Z(n2875) );
  OA31D0 U3137 ( .A1(n3226), .A2(n3218), .A3(n3227), .B(n2896), .Z(n3209) );
  OR2D0 U3138 ( .A1(n3228), .A2(n3229), .Z(n2896) );
  ND4D0 U3139 ( .A1(fifo_empty[7]), .A2(fifo_empty[6]), .A3(fifo_empty[5]), 
        .A4(fifo_empty[4]), .ZN(n3229) );
  ND4D0 U3140 ( .A1(fifo_empty[3]), .A2(fifo_empty[2]), .A3(fifo_empty[1]), 
        .A4(fifo_empty[0]), .ZN(n3228) );
  OAI31D0 U3141 ( .A1(n2930), .A2(n3055), .A3(n3230), .B(n3231), .ZN(n3227) );
  CKND2D0 U3142 ( .A1(n3107), .A2(n3001), .ZN(n2930) );
  ND4D0 U3143 ( .A1(n3232), .A2(n3216), .A3(n3215), .A4(n2969), .ZN(n3226) );
  CKND2D0 U3144 ( .A1(n3233), .A2(n3234), .ZN(n3225) );
  AOI221D0 U3145 ( .A1(n3212), .A2(n2938), .B1(n3213), .B2(n2939), .C(n3235), 
        .ZN(n3234) );
  OAI22D0 U3146 ( .A1(n2941), .A2(n3215), .B1(n2942), .B2(n3216), .ZN(n3235)
         );
  ND4D0 U3147 ( .A1(n3236), .A2(n3237), .A3(n2943), .A4(n3238), .ZN(n3216) );
  CKND0 U3148 ( .I(n3239), .ZN(n2942) );
  CKND2D0 U3149 ( .A1(n3080), .A2(n3236), .ZN(n3215) );
  CKND0 U3150 ( .I(n3232), .ZN(n3213) );
  CKND2D0 U3151 ( .A1(n2951), .A2(n3240), .ZN(n3232) );
  CKND0 U3152 ( .I(n3230), .ZN(n3212) );
  OAI31D0 U3153 ( .A1(n2950), .A2(n2948), .A3(n2952), .B(n3240), .ZN(n3230) );
  OA31D0 U3154 ( .A1(n2953), .A2(n2962), .A3(n2955), .B(n3241), .Z(n3240) );
  OR4D0 U3155 ( .A1(n3065), .A2(n3016), .A3(n3015), .A4(n3020), .Z(n2953) );
  ND4D0 U3156 ( .A1(n3068), .A2(n3066), .A3(n3242), .A4(n3067), .ZN(n2950) );
  NR2D0 U3157 ( .A1(n3010), .A2(n3012), .ZN(n3242) );
  AOI222D0 U3158 ( .A1(n3072), .A2(n2957), .B1(n3218), .B2(n2958), .C1(n3219), 
        .C2(n2959), .ZN(n3233) );
  CKND0 U3159 ( .I(n3231), .ZN(n3219) );
  CKND2D0 U3160 ( .A1(n2966), .A2(n3243), .ZN(n3231) );
  CKND0 U3161 ( .I(n3244), .ZN(n2966) );
  AN2D0 U3162 ( .A1(n2954), .A2(n3241), .Z(n3218) );
  OA211D0 U3163 ( .A1(n3245), .A2(n2964), .B(n3238), .C(n3236), .Z(n3241) );
  OA31D0 U3164 ( .A1(n2965), .A2(n2960), .A3(n2967), .B(n3243), .Z(n3236) );
  ND3D0 U3165 ( .A1(n2968), .A2(n2935), .A3(n2970), .ZN(n3243) );
  INR4D0 U3166 ( .A1(n3246), .B1(n3074), .B2(n3076), .B3(n3075), .ZN(n2970) );
  CKND0 U3167 ( .I(n3111), .ZN(n3075) );
  CKND0 U3168 ( .I(n3134), .ZN(n3076) );
  NR2D0 U3169 ( .A1(n2984), .A2(n3039), .ZN(n3246) );
  CKND0 U3170 ( .I(n3247), .ZN(n2960) );
  OR4D0 U3171 ( .A1(n3024), .A2(n3025), .A3(n3019), .A4(n3077), .Z(n2965) );
  CKND0 U3172 ( .I(n3248), .ZN(n3077) );
  ND3D0 U3173 ( .A1(n2971), .A2(n3173), .A3(n2973), .ZN(n3238) );
  INR4D0 U3174 ( .A1(n3249), .B1(n3056), .B2(n3002), .B3(n3083), .ZN(n2973) );
  CKND0 U3175 ( .I(n3206), .ZN(n3083) );
  NR2D0 U3176 ( .A1(n3084), .A2(n3082), .ZN(n3249) );
  CKND0 U3177 ( .I(n3137), .ZN(n3084) );
  CKND2D0 U3178 ( .A1(n3174), .A2(n3086), .ZN(n2964) );
  NR4D0 U3179 ( .A1(n3250), .A2(n3251), .A3(n3021), .A4(n3008), .ZN(n3174) );
  NR2D0 U3180 ( .A1(n3237), .A2(n2974), .ZN(n3245) );
  CKND2D0 U3181 ( .A1(n3252), .A2(n3253), .ZN(N3081) );
  AOI221D0 U3182 ( .A1(n3254), .A2(n2902), .B1(n3255), .B2(n2904), .C(n3256), 
        .ZN(n3253) );
  OAI22D0 U3183 ( .A1(n2906), .A2(n3257), .B1(n3258), .B2(n3259), .ZN(n3256)
         );
  CKND0 U3184 ( .I(n2913), .ZN(n3258) );
  ND4D0 U3185 ( .A1(n3260), .A2(n3261), .A3(n3262), .A4(n3263), .ZN(n2913) );
  NR3D0 U3186 ( .A1(n3264), .A2(n3265), .A3(n3266), .ZN(n3263) );
  AN4D0 U3187 ( .A1(n3267), .A2(n3268), .A3(n3269), .A4(n3270), .Z(n2906) );
  NR3D0 U3188 ( .A1(n3271), .A2(n3272), .A3(n3273), .ZN(n3270) );
  ND4D0 U3189 ( .A1(n3274), .A2(n3275), .A3(n3276), .A4(n3277), .ZN(n2904) );
  NR3D0 U3190 ( .A1(n3278), .A2(n3279), .A3(n3280), .ZN(n3277) );
  ND4D0 U3191 ( .A1(n3281), .A2(n3282), .A3(n3283), .A4(n3284), .ZN(n2902) );
  AOI222D0 U3192 ( .A1(n3074), .A2(n2911), .B1(n3285), .B2(n3217), .C1(n3286), 
        .C2(n2915), .ZN(n3252) );
  ND4D0 U3193 ( .A1(n3287), .A2(n3288), .A3(n3289), .A4(n3290), .ZN(n2915) );
  INR3D0 U3194 ( .A1(n3291), .B1(n3292), .B2(n3293), .ZN(n3290) );
  ND4D0 U3195 ( .A1(n3294), .A2(n3295), .A3(n3296), .A4(n3297), .ZN(n3217) );
  NR3D0 U3196 ( .A1(n3298), .A2(n3299), .A3(n3300), .ZN(n3297) );
  ND4D0 U3197 ( .A1(n3301), .A2(n3302), .A3(n3303), .A4(n3304), .ZN(n2911) );
  CKND2D0 U3198 ( .A1(n3305), .A2(n3306), .ZN(N3080) );
  AOI221D0 U3199 ( .A1(n3254), .A2(n2919), .B1(n3255), .B2(n2920), .C(n3307), 
        .ZN(n3306) );
  OAI22D0 U3200 ( .A1(n2922), .A2(n3257), .B1(n3308), .B2(n3259), .ZN(n3307)
         );
  CKND0 U3201 ( .I(n2925), .ZN(n3308) );
  ND4D0 U3202 ( .A1(n3309), .A2(n3261), .A3(n3310), .A4(n3311), .ZN(n2925) );
  AN4D0 U3203 ( .A1(n3312), .A2(n3268), .A3(n3313), .A4(n3314), .Z(n2922) );
  ND3D0 U3204 ( .A1(n3275), .A2(n3315), .A3(n3316), .ZN(n2920) );
  OAI211D0 U3205 ( .A1(n3317), .A2(n3318), .B(n3282), .C(n3281), .ZN(n2919) );
  NR2D0 U3206 ( .A1(n3319), .A2(n3320), .ZN(n3317) );
  AOI222D0 U3207 ( .A1(n3074), .A2(n2924), .B1(n3285), .B2(n3224), .C1(n3286), 
        .C2(n2926), .ZN(n3305) );
  ND4D0 U3208 ( .A1(n3321), .A2(n3288), .A3(n3322), .A4(n3323), .ZN(n2926) );
  ND4D0 U3209 ( .A1(n3324), .A2(n3295), .A3(n3325), .A4(n3326), .ZN(n3224) );
  ND3D0 U3210 ( .A1(n3302), .A2(n3327), .A3(n3328), .ZN(n2924) );
  CKND2D0 U3211 ( .A1(n3329), .A2(n3330), .ZN(N3079) );
  AOI221D0 U3212 ( .A1(n3254), .A2(n2938), .B1(n3255), .B2(n2939), .C(n3331), 
        .ZN(n3330) );
  OAI22D0 U3213 ( .A1(n2941), .A2(n3257), .B1(n3332), .B2(n3259), .ZN(n3331)
         );
  CKND2D0 U3214 ( .A1(n3065), .A2(n3333), .ZN(n3259) );
  NR3D0 U3215 ( .A1(n3334), .A2(n3335), .A3(n3336), .ZN(n3065) );
  CKND0 U3216 ( .I(n2958), .ZN(n3332) );
  IND4D0 U3217 ( .A1(n3264), .B1(n3309), .B2(n3337), .B3(n3338), .ZN(n2958) );
  INR2D0 U3218 ( .A1(n3339), .B1(n3340), .ZN(n3337) );
  AN3D0 U3219 ( .A1(n3260), .A2(n3341), .A3(n3262), .Z(n3309) );
  CKND2D0 U3220 ( .A1(n3082), .A2(n3342), .ZN(n3257) );
  CKND0 U3221 ( .I(n3136), .ZN(n3082) );
  ND3D0 U3222 ( .A1(n3343), .A2(n3344), .A3(n3345), .ZN(n3136) );
  IINR4D0 U3223 ( .A1(n3312), .A2(n3346), .B1(n3271), .B2(n3347), .ZN(n2941)
         );
  AN2D0 U3224 ( .A1(n3348), .A2(n3349), .Z(n3346) );
  AN3D0 U3225 ( .A1(n3267), .A2(n3350), .A3(n3269), .Z(n3312) );
  ND3D0 U3226 ( .A1(n3351), .A2(n3352), .A3(n3316), .ZN(n2939) );
  AN3D0 U3227 ( .A1(n3274), .A2(n3353), .A3(n3276), .Z(n3316) );
  INR2D0 U3228 ( .A1(n3354), .B1(n3068), .ZN(n3255) );
  ND3D0 U3229 ( .A1(n3355), .A2(n3356), .A3(n3357), .ZN(n3068) );
  IND4D0 U3230 ( .A1(n3320), .B1(n3281), .B2(n3283), .B3(n3358), .ZN(n2938) );
  AN4D0 U3231 ( .A1(n3359), .A2(n3360), .A3(n3361), .A4(n3362), .Z(n3281) );
  AN4D0 U3232 ( .A1(n3354), .A2(n3054), .A3(n3363), .A4(n3000), .Z(n3254) );
  CKND0 U3233 ( .I(n3107), .ZN(n3000) );
  OAI211D0 U3234 ( .A1(n3364), .A2(n3365), .B(n3362), .C(n3366), .ZN(n3107) );
  OAI21D0 U3235 ( .A1(n3367), .A2(n3368), .B(n3369), .ZN(n3362) );
  CKND0 U3236 ( .I(n3370), .ZN(n3368) );
  AOI31D0 U3237 ( .A1(n3371), .A2(n3372), .A3(n3373), .B(n3374), .ZN(n3367) );
  INR4D0 U3238 ( .A1(n3375), .B1(n3376), .B2(n3377), .B3(n3378), .ZN(n3364) );
  AOI21D0 U3239 ( .A1(n3379), .A2(n3380), .B(n3381), .ZN(n3378) );
  NR4D0 U3240 ( .A1(n3382), .A2(n3383), .A3(n3384), .A4(n3385), .ZN(n3380) );
  AOI211D0 U3241 ( .A1(n3386), .A2(n3387), .B(n3388), .C(n3389), .ZN(n3379) );
  ND4D0 U3242 ( .A1(n3390), .A2(n3391), .A3(n3392), .A4(n3393), .ZN(n3387) );
  CKND2D0 U3243 ( .A1(n3394), .A2(n3395), .ZN(n3376) );
  AOI31D0 U3244 ( .A1(n3066), .A2(n3067), .A3(n3204), .B(n3055), .ZN(n3363) );
  IND4D0 U3245 ( .A1(n3396), .B1(n3397), .B2(n3398), .B3(n3399), .ZN(n3055) );
  INR3D0 U3246 ( .A1(n3400), .B1(n3401), .B2(n3402), .ZN(n3399) );
  AOI211D0 U3247 ( .A1(n3403), .A2(n3404), .B(n3381), .C(n3365), .ZN(n3402) );
  NR4D0 U3248 ( .A1(n3405), .A2(n3406), .A3(n3383), .A4(n3385), .ZN(n3404) );
  AOI211D0 U3249 ( .A1(n3386), .A2(n3407), .B(n3408), .C(n3389), .ZN(n3403) );
  ND4D0 U3250 ( .A1(n3409), .A2(n3410), .A3(n3411), .A4(n3412), .ZN(n3407) );
  INR3D0 U3251 ( .A1(n3413), .B1(n3414), .B2(n3415), .ZN(n3412) );
  INR4D0 U3252 ( .A1(n3416), .B1(n2948), .B2(n2951), .B3(n3010), .ZN(n3204) );
  NR3D0 U3253 ( .A1(n3417), .A2(n3355), .A3(n3418), .ZN(n3010) );
  NR3D0 U3254 ( .A1(n3357), .A2(n3355), .A3(n3417), .ZN(n2951) );
  NR3D0 U3255 ( .A1(n3355), .A2(n3356), .A3(n3357), .ZN(n2948) );
  NR2D0 U3256 ( .A1(n3012), .A2(n2952), .ZN(n3416) );
  NR3D0 U3257 ( .A1(n3357), .A2(n3356), .A3(n3419), .ZN(n2952) );
  NR3D0 U3258 ( .A1(n3419), .A2(n3356), .A3(n3418), .ZN(n3012) );
  ND3D0 U3259 ( .A1(n3419), .A2(n3417), .A3(n3357), .ZN(n3067) );
  CKND0 U3260 ( .I(n3418), .ZN(n3357) );
  ND3D0 U3261 ( .A1(n3356), .A2(n3418), .A3(n3355), .ZN(n3066) );
  CKND0 U3262 ( .I(n3419), .ZN(n3355) );
  ND4D0 U3263 ( .A1(n3420), .A2(n3421), .A3(n3422), .A4(n3423), .ZN(n3419) );
  AOI211D0 U3264 ( .A1(n3424), .A2(n3425), .B(n3426), .C(n3427), .ZN(n3423) );
  OAI211D0 U3265 ( .A1(n3428), .A2(n3429), .B(n3430), .C(n3431), .ZN(n3425) );
  CKND0 U3266 ( .I(n3432), .ZN(n3430) );
  AOI211D0 U3267 ( .A1(n3433), .A2(n3434), .B(n3435), .C(n3436), .ZN(n3428) );
  OAI211D0 U3268 ( .A1(n3437), .A2(n3438), .B(n3439), .C(n3440), .ZN(n3435) );
  OAI211D0 U3269 ( .A1(n3441), .A2(n3442), .B(n3443), .C(n3444), .ZN(n3418) );
  NR2D0 U3270 ( .A1(n3445), .A2(n3446), .ZN(n3444) );
  OAI31D0 U3271 ( .A1(n3447), .A2(n3448), .A3(n3449), .B(n3424), .ZN(n3443) );
  AOI211D0 U3272 ( .A1(n3433), .A2(n3450), .B(n3451), .C(n3452), .ZN(n3441) );
  OAI21D0 U3273 ( .A1(n3453), .A2(n3438), .B(n3454), .ZN(n3451) );
  CKND0 U3274 ( .I(n3417), .ZN(n3356) );
  ND4D0 U3275 ( .A1(n3455), .A2(n3456), .A3(n3457), .A4(n3458), .ZN(n3417) );
  AN4D0 U3276 ( .A1(n3459), .A2(n3460), .A3(n3461), .A4(n3422), .Z(n3458) );
  INR2D0 U3277 ( .A1(n3462), .B1(n3427), .ZN(n3457) );
  OAI21D0 U3278 ( .A1(n3463), .A2(n3464), .B(n3424), .ZN(n3456) );
  OAI211D0 U3279 ( .A1(n3465), .A2(n3429), .B(n3466), .C(n3467), .ZN(n3464) );
  IINR4D0 U3280 ( .A1(n3468), .A2(n3469), .B1(n3470), .B2(n3471), .ZN(n3465)
         );
  OAI211D0 U3281 ( .A1(n3472), .A2(n3473), .B(n3474), .C(n3440), .ZN(n3470) );
  NR4D0 U3282 ( .A1(n3475), .A2(n3476), .A3(n3477), .A4(n3478), .ZN(n3472) );
  AOI31D0 U3283 ( .A1(n3479), .A2(n3480), .A3(n3481), .B(n3482), .ZN(n3478) );
  NR3D0 U3284 ( .A1(n3483), .A2(n3484), .A3(n3485), .ZN(n3481) );
  CKND0 U3285 ( .I(n3486), .ZN(n3479) );
  ND4D0 U3286 ( .A1(n3487), .A2(n3488), .A3(n3489), .A4(n3490), .ZN(n3463) );
  CKND0 U3287 ( .I(n3001), .ZN(n3054) );
  IND4D0 U3288 ( .A1(n3491), .B1(n3492), .B2(n3493), .B3(n3494), .ZN(n3001) );
  OA211D0 U3289 ( .A1(n3365), .A2(n3495), .B(n3496), .C(n3360), .Z(n3494) );
  AN4D0 U3290 ( .A1(n3375), .A2(n3497), .A3(n3498), .A4(n3499), .Z(n3495) );
  AOI211D0 U3291 ( .A1(n3500), .A2(n3501), .B(n3502), .C(n3503), .ZN(n3499) );
  ND4D0 U3292 ( .A1(n3504), .A2(n3505), .A3(n3506), .A4(n3507), .ZN(n3501) );
  NR4D0 U3293 ( .A1(n3405), .A2(n3406), .A3(n3382), .A4(n3384), .ZN(n3507) );
  CKND2D0 U3294 ( .A1(n3386), .A2(n3508), .ZN(n3505) );
  IND4D0 U3295 ( .A1(n3509), .B1(n3390), .B2(n3413), .B3(n3409), .ZN(n3508) );
  AN4D0 U3296 ( .A1(n3510), .A2(n3411), .A3(n3511), .A4(n3410), .Z(n3390) );
  NR2D0 U3297 ( .A1(n3512), .A2(n3513), .ZN(n3386) );
  OA21D0 U3298 ( .A1(n3016), .A2(n3123), .B(n3333), .Z(n3354) );
  OA211D0 U3299 ( .A1(n3250), .A2(n3514), .B(n3515), .C(n3342), .Z(n3333) );
  CKND0 U3300 ( .I(n3207), .ZN(n3514) );
  NR4D0 U3301 ( .A1(n3167), .A2(n3021), .A3(n3008), .A4(n2943), .ZN(n3207) );
  CKND0 U3302 ( .I(n2974), .ZN(n2943) );
  CKND2D0 U3303 ( .A1(n3516), .A2(n3517), .ZN(n2974) );
  NR3D0 U3304 ( .A1(n3516), .A2(n3518), .A3(n2945), .ZN(n3008) );
  NR3D0 U3305 ( .A1(n3516), .A2(n3237), .A3(n3517), .ZN(n3021) );
  CKND0 U3306 ( .I(n3086), .ZN(n3167) );
  ND3D0 U3307 ( .A1(n3516), .A2(n2945), .A3(n3518), .ZN(n3086) );
  CKND0 U3308 ( .I(n3085), .ZN(n3250) );
  NR2D0 U3309 ( .A1(n3129), .A2(n3117), .ZN(n3085) );
  NR3D0 U3310 ( .A1(n3518), .A2(n3237), .A3(n3516), .ZN(n3117) );
  NR3D0 U3311 ( .A1(n2945), .A2(n3519), .A3(n3517), .ZN(n3129) );
  OR4D0 U3312 ( .A1(n3520), .A2(n2955), .A3(n3015), .A4(n3020), .Z(n3123) );
  NR3D0 U3313 ( .A1(n3335), .A2(n3521), .A3(n3336), .ZN(n3020) );
  NR3D0 U3314 ( .A1(n3334), .A2(n3522), .A3(n3336), .ZN(n3015) );
  NR3D0 U3315 ( .A1(n3523), .A2(n3522), .A3(n3334), .ZN(n2955) );
  OR2D0 U3316 ( .A1(n2954), .A2(n2962), .Z(n3520) );
  NR3D0 U3317 ( .A1(n3522), .A2(n3521), .A3(n3523), .ZN(n2962) );
  NR3D0 U3318 ( .A1(n3523), .A2(n3521), .A3(n3335), .ZN(n2954) );
  OR2D0 U3319 ( .A1(n3128), .A2(n3124), .Z(n3016) );
  NR3D0 U3320 ( .A1(n3335), .A2(n3523), .A3(n3334), .ZN(n3124) );
  CKND0 U3321 ( .I(n3336), .ZN(n3523) );
  NR3D0 U3322 ( .A1(n3522), .A2(n3521), .A3(n3336), .ZN(n3128) );
  OAI221D0 U3323 ( .A1(n3524), .A2(n3525), .B1(n3526), .B2(n3527), .C(n3528), 
        .ZN(n3336) );
  NR2D0 U3324 ( .A1(n3529), .A2(n3530), .ZN(n3528) );
  AOI211D0 U3325 ( .A1(n3531), .A2(n3532), .B(n3533), .C(n3534), .ZN(n3524) );
  OAI21D0 U3326 ( .A1(n3535), .A2(n3536), .B(n3537), .ZN(n3533) );
  CKND0 U3327 ( .I(n3334), .ZN(n3521) );
  ND4D0 U3328 ( .A1(n3538), .A2(n3539), .A3(n3540), .A4(n3541), .ZN(n3334) );
  AOI211D0 U3329 ( .A1(n3542), .A2(n3543), .B(n3544), .C(n3545), .ZN(n3541) );
  ND4D0 U3330 ( .A1(n3546), .A2(n3547), .A3(n3548), .A4(n3549), .ZN(n3543) );
  AOI211D0 U3331 ( .A1(n3550), .A2(n3551), .B(n3552), .C(n3553), .ZN(n3549) );
  CKND0 U3332 ( .I(n3554), .ZN(n3553) );
  OAI211D0 U3333 ( .A1(n3555), .A2(n3556), .B(n3557), .C(n3558), .ZN(n3551) );
  AOI211D0 U3334 ( .A1(n3559), .A2(n3560), .B(n3561), .C(n3562), .ZN(n3558) );
  IND2D0 U3335 ( .A1(n3563), .B1(n3564), .ZN(n3560) );
  CKND0 U3336 ( .I(n3335), .ZN(n3522) );
  ND4D0 U3337 ( .A1(n3565), .A2(n3566), .A3(n3567), .A4(n3568), .ZN(n3335) );
  AN4D0 U3338 ( .A1(n3569), .A2(n3570), .A3(n3571), .A4(n3540), .Z(n3568) );
  INR2D0 U3339 ( .A1(n3572), .B1(n3545), .ZN(n3567) );
  OAI21D0 U3340 ( .A1(n3573), .A2(n3574), .B(n3542), .ZN(n3566) );
  OAI211D0 U3341 ( .A1(n3575), .A2(n3576), .B(n3577), .C(n3578), .ZN(n3574) );
  AN4D0 U3342 ( .A1(n3579), .A2(n3580), .A3(n3581), .A4(n3582), .Z(n3575) );
  OA211D0 U3343 ( .A1(n3583), .A2(n3536), .B(n3584), .C(n3585), .Z(n3579) );
  NR4D0 U3344 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3583) );
  AOI31D0 U3345 ( .A1(n3590), .A2(n3591), .A3(n3592), .B(n3593), .ZN(n3589) );
  NR3D0 U3346 ( .A1(n3594), .A2(n3595), .A3(n3596), .ZN(n3592) );
  ND4D0 U3347 ( .A1(n3554), .A2(n3548), .A3(n3597), .A4(n3598), .ZN(n3573) );
  AOI222D0 U3348 ( .A1(n3074), .A2(n2957), .B1(n3285), .B2(n3239), .C1(n3286), 
        .C2(n2959), .ZN(n3329) );
  ND4D0 U3349 ( .A1(n3321), .A2(n3291), .A3(n3599), .A4(n3600), .ZN(n2959) );
  INR2D0 U3350 ( .A1(n3601), .B1(n3602), .ZN(n3599) );
  AN3D0 U3351 ( .A1(n3287), .A2(n3603), .A3(n3289), .Z(n3321) );
  INR2D0 U3352 ( .A1(n3604), .B1(n3248), .ZN(n3286) );
  ND3D0 U3353 ( .A1(n3605), .A2(n3606), .A3(n3607), .ZN(n3248) );
  IND4D0 U3354 ( .A1(n3298), .B1(n3324), .B2(n3608), .B3(n3609), .ZN(n3239) );
  AN2D0 U3355 ( .A1(n3610), .A2(n3611), .Z(n3608) );
  AN3D0 U3356 ( .A1(n3294), .A2(n3612), .A3(n3296), .Z(n3324) );
  AN3D0 U3357 ( .A1(n3342), .A2(n3515), .A3(n3251), .Z(n3285) );
  CKND0 U3358 ( .I(n3087), .ZN(n3251) );
  ND3D0 U3359 ( .A1(n3237), .A2(n3519), .A3(n3518), .ZN(n3087) );
  CKND0 U3360 ( .I(n3517), .ZN(n3518) );
  ND4D0 U3361 ( .A1(n3613), .A2(n3614), .A3(n3615), .A4(n3616), .ZN(n3517) );
  AOI211D0 U3362 ( .A1(n3617), .A2(n3618), .B(n3619), .C(n3620), .ZN(n3616) );
  ND4D0 U3363 ( .A1(n3621), .A2(n3622), .A3(n3623), .A4(n3624), .ZN(n3618) );
  AOI211D0 U3364 ( .A1(n3625), .A2(n3626), .B(n3627), .C(n3628), .ZN(n3624) );
  CKND0 U3365 ( .I(n3629), .ZN(n3628) );
  IND4D0 U3366 ( .A1(n3630), .B1(n3631), .B2(n3632), .B3(n3633), .ZN(n3626) );
  AO31D0 U3367 ( .A1(n3634), .A2(n3635), .A3(n3636), .B(n3637), .Z(n3631) );
  OA21D0 U3368 ( .A1(n3638), .A2(n3639), .B(n3325), .Z(n3634) );
  CKND0 U3369 ( .I(n3516), .ZN(n3519) );
  IND3D0 U3370 ( .A1(n3640), .B1(n3641), .B2(n3642), .ZN(n3516) );
  OAI222D0 U3371 ( .A1(n3643), .A2(n3644), .B1(n3645), .B2(n3646), .C1(n3647), 
        .C2(n3648), .ZN(n3640) );
  NR2D0 U3372 ( .A1(n3649), .A2(n3650), .ZN(n3645) );
  AOI21D0 U3373 ( .A1(n3651), .A2(n3652), .B(n3653), .ZN(n3643) );
  CKND0 U3374 ( .I(n2945), .ZN(n3237) );
  ND4D0 U3375 ( .A1(n3654), .A2(n3655), .A3(n3656), .A4(n3657), .ZN(n2945) );
  AN4D0 U3376 ( .A1(n3658), .A2(n3659), .A3(n3660), .A4(n3615), .Z(n3657) );
  AOI21D0 U3377 ( .A1(n3617), .A2(n3661), .B(n3662), .ZN(n3656) );
  ND4D0 U3378 ( .A1(n3663), .A2(n3664), .A3(n3665), .A4(n3666), .ZN(n3661) );
  AN4D0 U3379 ( .A1(n3667), .A2(n3668), .A3(n3623), .A4(n3629), .Z(n3666) );
  OAI31D0 U3380 ( .A1(n3669), .A2(n3670), .A3(n3671), .B(n3625), .ZN(n3664) );
  AOI31D0 U3381 ( .A1(n3672), .A2(n3673), .A3(n3674), .B(n3637), .ZN(n3670) );
  AOI21D0 U3382 ( .A1(n3651), .A2(n3675), .B(n3676), .ZN(n3674) );
  OR4D0 U3383 ( .A1(n3677), .A2(n3678), .A3(n3679), .A4(n3680), .Z(n3675) );
  ND3D0 U3384 ( .A1(n3681), .A2(n3682), .A3(n3633), .ZN(n3669) );
  ND3D0 U3385 ( .A1(n3137), .A2(n3206), .A3(n3138), .ZN(n3515) );
  INR4D0 U3386 ( .A1(n3683), .B1(n3081), .B2(n3056), .B3(n3002), .ZN(n3138) );
  CKND0 U3387 ( .I(n3078), .ZN(n3002) );
  ND3D0 U3388 ( .A1(n3344), .A2(n3684), .A3(n3345), .ZN(n3078) );
  CKND0 U3389 ( .I(n3029), .ZN(n3056) );
  ND3D0 U3390 ( .A1(n3343), .A2(n3685), .A3(n3345), .ZN(n3029) );
  CKND0 U3391 ( .I(n2971), .ZN(n3081) );
  ND3D0 U3392 ( .A1(n3685), .A2(n3686), .A3(n3343), .ZN(n2971) );
  NR2D0 U3393 ( .A1(n3080), .A2(n2947), .ZN(n3683) );
  CKND0 U3394 ( .I(n3173), .ZN(n2947) );
  ND3D0 U3395 ( .A1(n3686), .A2(n3684), .A3(n3685), .ZN(n3173) );
  CKND0 U3396 ( .I(n2972), .ZN(n3080) );
  ND3D0 U3397 ( .A1(n3686), .A2(n3684), .A3(n3344), .ZN(n2972) );
  ND3D0 U3398 ( .A1(n3685), .A2(n3684), .A3(n3345), .ZN(n3206) );
  ND3D0 U3399 ( .A1(n3344), .A2(n3686), .A3(n3343), .ZN(n3137) );
  CKND0 U3400 ( .I(n3684), .ZN(n3343) );
  ND4D0 U3401 ( .A1(n3687), .A2(n3688), .A3(n3689), .A4(n3690), .ZN(n3684) );
  AOI211D0 U3402 ( .A1(n3691), .A2(n3692), .B(n3693), .C(n3694), .ZN(n3690) );
  ND4D0 U3403 ( .A1(n3695), .A2(n3696), .A3(n3697), .A4(n3698), .ZN(n3692) );
  AOI211D0 U3404 ( .A1(n3699), .A2(n3700), .B(n3701), .C(n3702), .ZN(n3698) );
  CKND0 U3405 ( .I(n3703), .ZN(n3702) );
  IND4D0 U3406 ( .A1(n3704), .B1(n3705), .B2(n3706), .B3(n3707), .ZN(n3700) );
  AO31D0 U3407 ( .A1(n3708), .A2(n3709), .A3(n3710), .B(n3711), .Z(n3705) );
  OA21D0 U3408 ( .A1(n3712), .A2(n3713), .B(n3313), .Z(n3708) );
  CKND0 U3409 ( .I(n3345), .ZN(n3686) );
  NR3D0 U3410 ( .A1(n3714), .A2(n3715), .A3(n3716), .ZN(n3345) );
  OAI222D0 U3411 ( .A1(n3717), .A2(n3718), .B1(n3719), .B2(n3720), .C1(n3721), 
        .C2(n3722), .ZN(n3716) );
  NR2D0 U3412 ( .A1(n3723), .A2(n3724), .ZN(n3719) );
  AOI21D0 U3413 ( .A1(n3725), .A2(n3726), .B(n3727), .ZN(n3717) );
  CKND0 U3414 ( .I(n3685), .ZN(n3344) );
  ND4D0 U3415 ( .A1(n3728), .A2(n3729), .A3(n3730), .A4(n3731), .ZN(n3685) );
  AN4D0 U3416 ( .A1(n3732), .A2(n3733), .A3(n3734), .A4(n3689), .Z(n3731) );
  AOI21D0 U3417 ( .A1(n3691), .A2(n3735), .B(n3736), .ZN(n3730) );
  ND4D0 U3418 ( .A1(n3737), .A2(n3738), .A3(n3739), .A4(n3740), .ZN(n3735) );
  AN4D0 U3419 ( .A1(n3741), .A2(n3742), .A3(n3697), .A4(n3703), .Z(n3740) );
  OAI31D0 U3420 ( .A1(n3743), .A2(n3744), .A3(n3745), .B(n3699), .ZN(n3738) );
  AOI31D0 U3421 ( .A1(n3746), .A2(n3747), .A3(n3748), .B(n3711), .ZN(n3744) );
  AOI21D0 U3422 ( .A1(n3725), .A2(n3749), .B(n3750), .ZN(n3748) );
  OR4D0 U3423 ( .A1(n3751), .A2(n3752), .A3(n3753), .A4(n3754), .Z(n3749) );
  ND3D0 U3424 ( .A1(n3755), .A2(n3756), .A3(n3707), .ZN(n3743) );
  OA21D0 U3425 ( .A1(n3025), .A2(n3131), .B(n3604), .Z(n3342) );
  ND3D0 U3426 ( .A1(n3134), .A2(n3111), .A3(n3135), .ZN(n3604) );
  INR4D0 U3427 ( .A1(n3757), .B1(n2910), .B2(n3072), .B3(n2984), .ZN(n3135) );
  CKND0 U3428 ( .I(n2995), .ZN(n2984) );
  ND3D0 U3429 ( .A1(n3758), .A2(n3759), .A3(n3760), .ZN(n2995) );
  CKND0 U3430 ( .I(n2969), .ZN(n3072) );
  ND3D0 U3431 ( .A1(n3761), .A2(n3759), .A3(n3758), .ZN(n2969) );
  CKND0 U3432 ( .I(n2935), .ZN(n2910) );
  ND3D0 U3433 ( .A1(n3761), .A2(n3759), .A3(n3762), .ZN(n2935) );
  NR2D0 U3434 ( .A1(n3039), .A2(n3073), .ZN(n3757) );
  CKND0 U3435 ( .I(n2968), .ZN(n3073) );
  ND3D0 U3436 ( .A1(n3762), .A2(n3761), .A3(n3763), .ZN(n2968) );
  CKND0 U3437 ( .I(n3027), .ZN(n3039) );
  ND3D0 U3438 ( .A1(n3763), .A2(n3762), .A3(n3760), .ZN(n3027) );
  ND3D0 U3439 ( .A1(n3762), .A2(n3759), .A3(n3760), .ZN(n3111) );
  ND3D0 U3440 ( .A1(n3758), .A2(n3761), .A3(n3763), .ZN(n3134) );
  IND4D0 U3441 ( .A1(n3019), .B1(n3247), .B2(n3244), .B3(n3764), .ZN(n3131) );
  NR2D0 U3442 ( .A1(n3024), .A2(n2967), .ZN(n3764) );
  NR3D0 U3443 ( .A1(n3607), .A2(n3606), .A3(n3765), .ZN(n2967) );
  NR3D0 U3444 ( .A1(n3765), .A2(n3606), .A3(n3766), .ZN(n3024) );
  ND3D0 U3445 ( .A1(n3766), .A2(n3765), .A3(n3606), .ZN(n3244) );
  ND3D0 U3446 ( .A1(n3767), .A2(n3765), .A3(n3766), .ZN(n3247) );
  NR3D0 U3447 ( .A1(n3767), .A2(n3605), .A3(n3766), .ZN(n3019) );
  OR2D0 U3448 ( .A1(n3126), .A2(n3132), .Z(n3025) );
  NR3D0 U3449 ( .A1(n3767), .A2(n3607), .A3(n3765), .ZN(n3132) );
  CKND0 U3450 ( .I(n3605), .ZN(n3765) );
  CKND0 U3451 ( .I(n3766), .ZN(n3607) );
  NR3D0 U3452 ( .A1(n3606), .A2(n3605), .A3(n3766), .ZN(n3126) );
  OAI211D0 U3453 ( .A1(n3768), .A2(n3769), .B(n3289), .C(n3770), .ZN(n3766) );
  AOI21D0 U3454 ( .A1(n3771), .A2(n3772), .B(n3773), .ZN(n3770) );
  CKND2D0 U3455 ( .A1(n3774), .A2(n3775), .ZN(n3772) );
  AOI211D0 U3456 ( .A1(n3776), .A2(n3777), .B(n3778), .C(n3779), .ZN(n3768) );
  OAI211D0 U3457 ( .A1(n3780), .A2(n3781), .B(n3782), .C(n3783), .ZN(n3777) );
  AOI21D0 U3458 ( .A1(n3784), .A2(n3785), .B(n3786), .ZN(n3783) );
  INR3D0 U3459 ( .A1(n3787), .B1(n3788), .B2(n3789), .ZN(n3605) );
  AOI211D0 U3460 ( .A1(n3790), .A2(n3791), .B(n3792), .C(n3793), .ZN(n3787) );
  ND4D0 U3461 ( .A1(n3794), .A2(n3795), .A3(n3796), .A4(n3797), .ZN(n3791) );
  AOI211D0 U3462 ( .A1(n3776), .A2(n3798), .B(n3799), .C(n3800), .ZN(n3797) );
  IND4D0 U3463 ( .A1(n3801), .B1(n3802), .B2(n3803), .B3(n3804), .ZN(n3798) );
  OAI31D0 U3464 ( .A1(n3805), .A2(n3806), .A3(n3807), .B(n3808), .ZN(n3802) );
  OAI21D0 U3465 ( .A1(n3809), .A2(n3810), .B(n3811), .ZN(n3805) );
  CKND0 U3466 ( .I(n3767), .ZN(n3606) );
  ND4D0 U3467 ( .A1(n3812), .A2(n3813), .A3(n3814), .A4(n3815), .ZN(n3767) );
  NR4D0 U3468 ( .A1(n3816), .A2(n3817), .A3(n3793), .A4(n3818), .ZN(n3815) );
  CKND2D0 U3469 ( .A1(n3790), .A2(n3819), .ZN(n3813) );
  ND4D0 U3470 ( .A1(n3820), .A2(n3821), .A3(n3822), .A4(n3823), .ZN(n3819) );
  AN4D0 U3471 ( .A1(n3824), .A2(n3825), .A3(n3796), .A4(n3826), .Z(n3823) );
  OAI31D0 U3472 ( .A1(n3827), .A2(n3828), .A3(n3829), .B(n3776), .ZN(n3821) );
  AOI31D0 U3473 ( .A1(n3830), .A2(n3831), .A3(n3832), .B(n3781), .ZN(n3828) );
  OA21D0 U3474 ( .A1(n3810), .A2(n3833), .B(n3834), .Z(n3832) );
  AN4D0 U3475 ( .A1(n3835), .A2(n3836), .A3(n3837), .A4(n3838), .Z(n3833) );
  ND3D0 U3476 ( .A1(n3804), .A2(n3839), .A3(n3840), .ZN(n3827) );
  CKND0 U3477 ( .I(n3769), .ZN(n3790) );
  ND3D0 U3478 ( .A1(n3303), .A2(n3841), .A3(n3328), .ZN(n2957) );
  AN2D0 U3479 ( .A1(n3301), .A2(n3842), .Z(n3328) );
  AN4D0 U3480 ( .A1(n3843), .A2(n3844), .A3(n3845), .A4(n3846), .Z(n3301) );
  INR2D0 U3481 ( .A1(n3847), .B1(n3848), .ZN(n3845) );
  CKND0 U3482 ( .I(n3133), .ZN(n3074) );
  ND3D0 U3483 ( .A1(n3763), .A2(n3758), .A3(n3760), .ZN(n3133) );
  CKND0 U3484 ( .I(n3761), .ZN(n3760) );
  OAI221D0 U3485 ( .A1(n3849), .A2(n3850), .B1(n3851), .B2(n3844), .C(n3843), 
        .ZN(n3761) );
  AN3D0 U3486 ( .A1(n3852), .A2(n3853), .A3(n3854), .Z(n3843) );
  AOI221D0 U3487 ( .A1(n3855), .A2(n3856), .B1(n3857), .B2(n3858), .C(n3859), 
        .ZN(n3849) );
  OAI221D0 U3488 ( .A1(n3860), .A2(n3861), .B1(n3862), .B2(n3863), .C(n3864), 
        .ZN(n3856) );
  AOI221D0 U3489 ( .A1(n3865), .A2(n3866), .B1(n3867), .B2(n3865), .C(n3868), 
        .ZN(n3860) );
  CKND0 U3490 ( .I(n3869), .ZN(n3868) );
  OAI221D0 U3491 ( .A1(n3870), .A2(n3871), .B1(n3872), .B2(n3873), .C(n3874), 
        .ZN(n3866) );
  AOI221D0 U3492 ( .A1(n3875), .A2(n3876), .B1(n3877), .B2(n3878), .C(n3879), 
        .ZN(n3870) );
  OAI221D0 U3493 ( .A1(n3880), .A2(n3881), .B1(n3882), .B2(n3883), .C(n3884), 
        .ZN(n3876) );
  AOI31D0 U3494 ( .A1(n3885), .A2(n3886), .A3(n3887), .B(n3888), .ZN(n3880) );
  CKND0 U3495 ( .I(n3762), .ZN(n3758) );
  OAI211D0 U3496 ( .A1(n3889), .A2(n3850), .B(n3890), .C(n3891), .ZN(n3762) );
  INR2D0 U3497 ( .A1(n3854), .B1(n3892), .ZN(n3891) );
  NR4D0 U3498 ( .A1(n3893), .A2(n3894), .A3(n3895), .A4(n3896), .ZN(n3892) );
  ND4D0 U3499 ( .A1(n3897), .A2(n3898), .A3(n3899), .A4(n3900), .ZN(n3854) );
  NR2D0 U3500 ( .A1(n3901), .A2(n3372), .ZN(n3899) );
  AOI221D0 U3501 ( .A1(n3902), .A2(n3903), .B1(n3855), .B2(n3904), .C(n3905), 
        .ZN(n3889) );
  OAI211D0 U3502 ( .A1(n3906), .A2(n3861), .B(n3907), .C(n3908), .ZN(n3904) );
  AOI21D0 U3503 ( .A1(n3909), .A2(n3910), .B(n3911), .ZN(n3908) );
  CKND0 U3504 ( .I(n3912), .ZN(n3911) );
  CKND0 U3505 ( .I(n3913), .ZN(n3907) );
  AOI221D0 U3506 ( .A1(n3865), .A2(n3914), .B1(n3915), .B2(n3916), .C(n3917), 
        .ZN(n3906) );
  OAI211D0 U3507 ( .A1(n3918), .A2(n3871), .B(n3919), .C(n3920), .ZN(n3914) );
  AOI21D0 U3508 ( .A1(n3921), .A2(n3922), .B(n3923), .ZN(n3920) );
  AOI221D0 U3509 ( .A1(n3875), .A2(n3924), .B1(n3925), .B2(n3926), .C(n3927), 
        .ZN(n3918) );
  CKND0 U3510 ( .I(n3928), .ZN(n3927) );
  OAI211D0 U3511 ( .A1(n3929), .A2(n3930), .B(n3931), .C(n3932), .ZN(n3924) );
  AOI21D0 U3512 ( .A1(n3933), .A2(n3934), .B(n3935), .ZN(n3932) );
  CKND0 U3513 ( .I(n3936), .ZN(n3935) );
  OAI21D0 U3514 ( .A1(n3937), .A2(n3895), .B(n3938), .ZN(n3934) );
  CKND0 U3515 ( .I(n3939), .ZN(n3931) );
  CKND0 U3516 ( .I(n3940), .ZN(n3929) );
  CKND0 U3517 ( .I(n3759), .ZN(n3763) );
  OAI211D0 U3518 ( .A1(n3848), .A2(n3846), .B(n3890), .C(n3941), .ZN(n3759) );
  AOI21D0 U3519 ( .A1(n3942), .A2(n3943), .B(n3944), .ZN(n3941) );
  CKND0 U3520 ( .I(n3853), .ZN(n3944) );
  ND4D0 U3521 ( .A1(n3942), .A2(n3898), .A3(n3945), .A4(n3946), .ZN(n3853) );
  OAI221D0 U3522 ( .A1(n3947), .A2(n3948), .B1(n3949), .B2(n3950), .C(n3951), 
        .ZN(n3943) );
  AOI211D0 U3523 ( .A1(n3952), .A2(n3953), .B(n3954), .C(n3913), .ZN(n3947) );
  OAI211D0 U3524 ( .A1(n3955), .A2(n3861), .B(n3956), .C(n3957), .ZN(n3913) );
  ND4D0 U3525 ( .A1(n3953), .A2(n3958), .A3(n3959), .A4(n3960), .ZN(n3956) );
  NR2D0 U3526 ( .A1(n3952), .A2(n3961), .ZN(n3959) );
  NR2D0 U3527 ( .A1(n3962), .A2(n3963), .ZN(n3955) );
  OAI221D0 U3528 ( .A1(n3964), .A2(n3965), .B1(n3966), .B2(n3861), .C(n3967), 
        .ZN(n3954) );
  AOI221D0 U3529 ( .A1(n3968), .A2(n3969), .B1(n3865), .B2(n3970), .C(n3971), 
        .ZN(n3966) );
  OAI211D0 U3530 ( .A1(n3972), .A2(n3973), .B(n3919), .C(n3974), .ZN(n3970) );
  AOI21D0 U3531 ( .A1(n3975), .A2(n3976), .B(n3977), .ZN(n3974) );
  OAI22D0 U3532 ( .A1(n3978), .A2(n3979), .B1(n3980), .B2(n3981), .ZN(n3976)
         );
  AOI211D0 U3533 ( .A1(n3982), .A2(n3983), .B(n3984), .C(n3939), .ZN(n3980) );
  OAI211D0 U3534 ( .A1(n3985), .A2(n3881), .B(n3986), .C(n3987), .ZN(n3939) );
  AN2D0 U3535 ( .A1(n3988), .A2(n3989), .Z(n3985) );
  OAI221D0 U3536 ( .A1(n3990), .A2(n3991), .B1(n3992), .B2(n3881), .C(n3993), 
        .ZN(n3984) );
  CKND0 U3537 ( .I(n3933), .ZN(n3881) );
  OA21D0 U3538 ( .A1(n3994), .A2(n3995), .B(n3996), .Z(n3992) );
  CKND2D0 U3539 ( .A1(n3930), .A2(n3940), .ZN(n3991) );
  OA211D0 U3540 ( .A1(n3997), .A2(n3871), .B(n3998), .C(n3999), .Z(n3919) );
  ND4D0 U3541 ( .A1(n4000), .A2(n4001), .A3(n4002), .A4(n3960), .ZN(n3998) );
  NR2D0 U3542 ( .A1(n4003), .A2(n4004), .ZN(n4002) );
  INR2D0 U3543 ( .A1(n4005), .B1(n4006), .ZN(n3997) );
  CKND0 U3544 ( .I(n4000), .ZN(n3972) );
  AN3D0 U3545 ( .A1(n3847), .A2(n3852), .A3(n4007), .Z(n3890) );
  ND3D0 U3546 ( .A1(n3942), .A2(n3898), .A3(n4008), .ZN(n3852) );
  AOI211D0 U3547 ( .A1(n3945), .A2(n3946), .B(n4009), .C(n3373), .ZN(n4008) );
  CKND0 U3548 ( .I(n3850), .ZN(n3942) );
  CKND2D0 U3549 ( .A1(n4010), .A2(n3897), .ZN(n3850) );
  CKND0 U3550 ( .I(n3851), .ZN(n3897) );
  OAI31D0 U3551 ( .A1(n3896), .A2(n4011), .A3(n4012), .B(n4013), .ZN(n3851) );
  AOI31D0 U3552 ( .A1(n3900), .A2(n4014), .A3(n3898), .B(n3901), .ZN(n4010) );
  CKND0 U3553 ( .I(n3844), .ZN(n3901) );
  ND3D0 U3554 ( .A1(n4015), .A2(n4016), .A3(n3898), .ZN(n3844) );
  IND4D0 U3555 ( .A1(n4011), .B1(n4013), .B2(n3898), .B3(n3960), .ZN(n3847) );
  NR2D0 U3556 ( .A1(n3848), .A2(n4017), .ZN(n4013) );
  CKND0 U3557 ( .I(n3846), .ZN(n4017) );
  ND3D0 U3558 ( .A1(n4018), .A2(n4019), .A3(n3898), .ZN(n3846) );
  CKND0 U3559 ( .I(n3896), .ZN(n3898) );
  INR2D0 U3560 ( .A1(n4020), .B1(n3896), .ZN(n3848) );
  CKND2D0 U3561 ( .A1(n3302), .A2(n4021), .ZN(n3896) );
  IINR4D0 U3562 ( .A1(n4007), .A2(n4022), .B1(n3859), .B2(n3857), .ZN(n3302)
         );
  OAI31D0 U3563 ( .A1(n3965), .A2(n3964), .A3(n3948), .B(n4023), .ZN(n3859) );
  CKND0 U3564 ( .I(n3905), .ZN(n4023) );
  OAI31D0 U3565 ( .A1(n4024), .A2(n3964), .A3(n4025), .B(n3951), .ZN(n3905) );
  ND4D0 U3566 ( .A1(n3855), .A2(n4021), .A3(n4026), .A4(n4027), .ZN(n3951) );
  AN2D0 U3567 ( .A1(n4028), .A2(n3965), .Z(n4026) );
  CKND0 U3568 ( .I(n3948), .ZN(n3855) );
  ND3D0 U3569 ( .A1(n4029), .A2(n4030), .A3(n3900), .ZN(n4024) );
  CKND2D0 U3570 ( .A1(n4031), .A2(n3858), .ZN(n3948) );
  CKND0 U3571 ( .I(n4025), .ZN(n3858) );
  CKND2D0 U3572 ( .A1(n4022), .A2(n4032), .ZN(n4025) );
  AOI31D0 U3573 ( .A1(n3900), .A2(n4029), .A3(n4021), .B(n3857), .ZN(n4031) );
  CKND0 U3574 ( .I(n4030), .ZN(n3857) );
  ND3D0 U3575 ( .A1(n4015), .A2(n4033), .A3(n4021), .ZN(n4030) );
  CKND2D0 U3576 ( .A1(n3945), .A2(n4034), .ZN(n3965) );
  IND2D0 U3577 ( .A1(n4032), .B1(n4022), .ZN(n4007) );
  INR2D0 U3578 ( .A1(n3950), .B1(n3949), .ZN(n4022) );
  AO21D0 U3579 ( .A1(n4035), .A2(n4021), .B(n3902), .Z(n3949) );
  NR3D0 U3580 ( .A1(n3895), .A2(n4036), .A3(n3964), .ZN(n3902) );
  ND3D0 U3581 ( .A1(n4018), .A2(n4037), .A3(n4021), .ZN(n3950) );
  ND3D0 U3582 ( .A1(n3960), .A2(n4038), .A3(n4021), .ZN(n4032) );
  CKND0 U3583 ( .I(n3964), .ZN(n4021) );
  CKND2D0 U3584 ( .A1(n3303), .A2(n3958), .ZN(n3964) );
  AN2D0 U3585 ( .A1(n3864), .A2(n4039), .Z(n3303) );
  AN3D0 U3586 ( .A1(n3912), .A2(n3967), .A3(n3957), .Z(n3864) );
  ND3D0 U3587 ( .A1(n4040), .A2(n3958), .A3(n4041), .ZN(n3957) );
  AOI211D0 U3588 ( .A1(n3945), .A2(n4042), .B(n4009), .C(n4043), .ZN(n4041) );
  ND4D0 U3589 ( .A1(n4040), .A2(n3958), .A3(n3945), .A4(n4042), .ZN(n3967) );
  CKND0 U3590 ( .I(n3861), .ZN(n4040) );
  OAI31D0 U3591 ( .A1(n4044), .A2(n4045), .A3(n4046), .B(n4039), .ZN(n3861) );
  ND4D0 U3592 ( .A1(n4039), .A2(n3958), .A3(n3900), .A4(n4047), .ZN(n3912) );
  INR2D0 U3593 ( .A1(n3863), .B1(n3862), .ZN(n4039) );
  CKND2D0 U3594 ( .A1(n4048), .A2(n3953), .ZN(n3862) );
  AOI21D0 U3595 ( .A1(n4049), .A2(n3958), .B(n3909), .ZN(n3953) );
  NR3D0 U3596 ( .A1(n3895), .A2(n4050), .A3(n4044), .ZN(n3909) );
  AOI31D0 U3597 ( .A1(n3960), .A2(n4051), .A3(n3958), .B(n3952), .ZN(n4048) );
  AN3D0 U3598 ( .A1(n4018), .A2(n4052), .A3(n3958), .Z(n3952) );
  ND3D0 U3599 ( .A1(n4015), .A2(n4053), .A3(n3958), .ZN(n3863) );
  CKND0 U3600 ( .I(n4044), .ZN(n3958) );
  CKND2D0 U3601 ( .A1(n3304), .A2(n4054), .ZN(n4044) );
  AN4D0 U3602 ( .A1(n3869), .A2(n3969), .A3(n4055), .A4(n4056), .Z(n3304) );
  NR2D0 U3603 ( .A1(n3963), .A2(n3968), .ZN(n4055) );
  INR3D0 U3604 ( .A1(n3969), .B1(n4057), .B2(n3968), .ZN(n3963) );
  CKND0 U3605 ( .I(n4058), .ZN(n3968) );
  NR3D0 U3606 ( .A1(n3971), .A2(n3917), .A3(n3962), .ZN(n3869) );
  AN4D0 U3607 ( .A1(n4059), .A2(n4027), .A3(n4060), .A4(n4061), .Z(n3962) );
  CKND2D0 U3608 ( .A1(n3945), .A2(n4062), .ZN(n4061) );
  INR4D0 U3609 ( .A1(n3865), .B1(n4063), .B2(n4064), .B3(n3867), .ZN(n3917) );
  CKND0 U3610 ( .I(n4056), .ZN(n3867) );
  AN3D0 U3611 ( .A1(n3945), .A2(n4062), .A3(n4059), .Z(n3971) );
  AN4D0 U3612 ( .A1(n3865), .A2(n4054), .A3(n4056), .A4(n4063), .Z(n4059) );
  CKND2D0 U3613 ( .A1(n3900), .A2(n4065), .ZN(n4063) );
  ND3D0 U3614 ( .A1(n4015), .A2(n4066), .A3(n4054), .ZN(n4056) );
  AN3D0 U3615 ( .A1(n4057), .A2(n4058), .A3(n3969), .Z(n3865) );
  AOI21D0 U3616 ( .A1(n4067), .A2(n4054), .B(n3915), .ZN(n3969) );
  NR3D0 U3617 ( .A1(n3895), .A2(n4068), .A3(n4064), .ZN(n3915) );
  ND3D0 U3618 ( .A1(n4018), .A2(n4069), .A3(n4054), .ZN(n4058) );
  ND3D0 U3619 ( .A1(n3960), .A2(n4070), .A3(n4054), .ZN(n4057) );
  CKND0 U3620 ( .I(n4064), .ZN(n4054) );
  CKND2D0 U3621 ( .A1(n3842), .A2(n4001), .ZN(n4064) );
  AN2D0 U3622 ( .A1(n3874), .A2(n4071), .Z(n3842) );
  INR3D0 U3623 ( .A1(n3999), .B1(n3923), .B2(n3977), .ZN(n3874) );
  INR4D0 U3624 ( .A1(n3945), .B1(n3871), .B2(n4072), .B3(n4073), .ZN(n3977) );
  INR4D0 U3625 ( .A1(n4071), .B1(n4072), .B2(n4046), .B3(n4074), .ZN(n3923) );
  ND3D0 U3626 ( .A1(n3975), .A2(n4001), .A3(n4075), .ZN(n3999) );
  AOI211D0 U3627 ( .A1(n3945), .A2(n4076), .B(n4009), .C(n4077), .ZN(n4075) );
  CKND0 U3628 ( .I(n3871), .ZN(n3975) );
  OAI31D0 U3629 ( .A1(n4072), .A2(n4074), .A3(n4046), .B(n4071), .ZN(n3871) );
  INR2D0 U3630 ( .A1(n3873), .B1(n3872), .ZN(n4071) );
  CKND2D0 U3631 ( .A1(n4078), .A2(n4000), .ZN(n3872) );
  AOI21D0 U3632 ( .A1(n4079), .A2(n4001), .B(n3921), .ZN(n4000) );
  NR3D0 U3633 ( .A1(n3895), .A2(n4080), .A3(n4072), .ZN(n3921) );
  AOI31D0 U3634 ( .A1(n3960), .A2(n4081), .A3(n4001), .B(n4003), .ZN(n4078) );
  CKND0 U3635 ( .I(n3973), .ZN(n4003) );
  ND3D0 U3636 ( .A1(n4018), .A2(n4082), .A3(n4001), .ZN(n3973) );
  ND3D0 U3637 ( .A1(n4015), .A2(n4083), .A3(n4001), .ZN(n3873) );
  CKND0 U3638 ( .I(n4072), .ZN(n4001) );
  CKND2D0 U3639 ( .A1(n3327), .A2(n3983), .ZN(n4072) );
  INR4D0 U3640 ( .A1(n4084), .B1(n3879), .B2(n3978), .B3(n3877), .ZN(n3327) );
  OAI211D0 U3641 ( .A1(n4085), .A2(n4086), .B(n4005), .C(n3928), .ZN(n3879) );
  ND4D0 U3642 ( .A1(n4087), .A2(n4088), .A3(n3900), .A4(n4089), .ZN(n3928) );
  INR2D0 U3643 ( .A1(n3878), .B1(n4090), .ZN(n4089) );
  ND4D0 U3644 ( .A1(n3875), .A2(n3983), .A3(n4091), .A4(n4027), .ZN(n4005) );
  NR2D0 U3645 ( .A1(n3982), .A2(n4092), .ZN(n4091) );
  CKND0 U3646 ( .I(n4085), .ZN(n3982) );
  CKND2D0 U3647 ( .A1(n3875), .A2(n3983), .ZN(n4086) );
  CKND0 U3648 ( .I(n3981), .ZN(n3875) );
  CKND2D0 U3649 ( .A1(n4093), .A2(n3878), .ZN(n3981) );
  INR3D0 U3650 ( .A1(n4094), .B1(n4095), .B2(n3978), .ZN(n3878) );
  AOI31D0 U3651 ( .A1(n3900), .A2(n4087), .A3(n3983), .B(n3877), .ZN(n4093) );
  CKND0 U3652 ( .I(n4088), .ZN(n3877) );
  ND3D0 U3653 ( .A1(n4015), .A2(n4096), .A3(n3983), .ZN(n4088) );
  CKND2D0 U3654 ( .A1(n3945), .A2(n4097), .ZN(n4085) );
  NR2D0 U3655 ( .A1(n4006), .A2(n4095), .ZN(n4084) );
  NR3D0 U3656 ( .A1(n4094), .A2(n4095), .A3(n3978), .ZN(n4006) );
  AO21D0 U3657 ( .A1(n4098), .A2(n3983), .B(n3925), .Z(n3978) );
  NR3D0 U3658 ( .A1(n3895), .A2(n4099), .A3(n4090), .ZN(n3925) );
  CKND0 U3659 ( .I(n3979), .ZN(n4095) );
  ND3D0 U3660 ( .A1(n4018), .A2(n4100), .A3(n3983), .ZN(n3979) );
  ND3D0 U3661 ( .A1(n3960), .A2(n4101), .A3(n3983), .ZN(n4094) );
  CKND0 U3662 ( .I(n4090), .ZN(n3983) );
  CKND2D0 U3663 ( .A1(n3841), .A2(n4102), .ZN(n4090) );
  AN4D0 U3664 ( .A1(n3884), .A2(n4103), .A3(n3986), .A4(n3883), .Z(n3841) );
  ND4D0 U3665 ( .A1(n4103), .A2(n4102), .A3(n3960), .A4(n4104), .ZN(n3986) );
  AN3D0 U3666 ( .A1(n3993), .A2(n3936), .A3(n3987), .Z(n3884) );
  ND3D0 U3667 ( .A1(n3933), .A2(n4102), .A3(n4105), .ZN(n3987) );
  AOI211D0 U3668 ( .A1(n3945), .A2(n4106), .B(n4009), .C(n4107), .ZN(n4105) );
  IND3D0 U3669 ( .A1(n3882), .B1(n3883), .B2(n4108), .ZN(n3936) );
  ND4D0 U3670 ( .A1(n3933), .A2(n4102), .A3(n3945), .A4(n4106), .ZN(n3993) );
  INR3D0 U3671 ( .A1(n3883), .B1(n4108), .B2(n3882), .ZN(n3933) );
  OAI31D0 U3672 ( .A1(n4109), .A2(n4110), .A3(n4012), .B(n4103), .ZN(n3882) );
  AN3D0 U3673 ( .A1(n3990), .A2(n3940), .A3(n3930), .Z(n4103) );
  IND3D0 U3674 ( .A1(n3895), .B1(n4111), .B2(n4102), .ZN(n3930) );
  CKND2D0 U3675 ( .A1(n4102), .A2(n4112), .ZN(n3940) );
  ND3D0 U3676 ( .A1(n4018), .A2(n4113), .A3(n4102), .ZN(n3990) );
  NR3D0 U3677 ( .A1(n4046), .A2(n4114), .A3(n4109), .ZN(n4108) );
  ND3D0 U3678 ( .A1(n4015), .A2(n4115), .A3(n4102), .ZN(n3883) );
  CKND0 U3679 ( .I(n4109), .ZN(n4102) );
  IND4D0 U3680 ( .A1(n3888), .B1(n3885), .B2(n3988), .B3(n4116), .ZN(n4109) );
  CKND2D0 U3681 ( .A1(n3885), .A2(n4117), .ZN(n3988) );
  ND3D0 U3682 ( .A1(n3996), .A2(n3938), .A3(n3989), .ZN(n3888) );
  ND4D0 U3683 ( .A1(n4027), .A2(n4118), .A3(n4119), .A4(n4120), .ZN(n3989) );
  CKND2D0 U3684 ( .A1(n3945), .A2(n4121), .ZN(n4120) );
  CKND0 U3685 ( .I(n4009), .ZN(n4027) );
  OAI221D0 U3686 ( .A1(n4122), .A2(n4123), .B1(n4124), .B2(n3769), .C(n3812), 
        .ZN(n4009) );
  CKND0 U3687 ( .I(n4125), .ZN(n3812) );
  AOI221D0 U3688 ( .A1(n4126), .A2(n4127), .B1(n3776), .B2(n4128), .C(n4129), 
        .ZN(n4124) );
  OAI221D0 U3689 ( .A1(n3838), .A2(n4130), .B1(n4123), .B2(n4131), .C(n4132), 
        .ZN(n4128) );
  CKND0 U3690 ( .I(n3829), .ZN(n4132) );
  NR4D0 U3691 ( .A1(n4133), .A2(n4134), .A3(n4135), .A4(n4136), .ZN(n4131) );
  IND3D0 U3692 ( .A1(n4137), .B1(n3837), .B2(n4138), .ZN(n4133) );
  IND3D0 U3693 ( .A1(n4139), .B1(n4140), .B2(n3822), .ZN(n4127) );
  NR3D0 U3694 ( .A1(n4141), .A2(n4142), .A3(n4143), .ZN(n4122) );
  ND3D0 U3695 ( .A1(n3900), .A2(n4144), .A3(n4145), .ZN(n3938) );
  CKND0 U3696 ( .I(n4046), .ZN(n3900) );
  ND3D0 U3697 ( .A1(n4118), .A2(n4121), .A3(n3945), .ZN(n3996) );
  OA21D0 U3698 ( .A1(n4146), .A2(n4046), .B(n4145), .Z(n4118) );
  INR3D0 U3699 ( .A1(n3885), .B1(n4117), .B2(n3887), .ZN(n4145) );
  CKND0 U3700 ( .I(n4116), .ZN(n3887) );
  CKND2D0 U3701 ( .A1(n4015), .A2(n4147), .ZN(n4116) );
  CKND0 U3702 ( .I(n3886), .ZN(n4117) );
  CKND2D0 U3703 ( .A1(n3960), .A2(n4148), .ZN(n3886) );
  INR2D0 U3704 ( .A1(n3994), .B1(n3995), .ZN(n3885) );
  OAI21D0 U3705 ( .A1(n4149), .A2(n3895), .B(n4150), .ZN(n3995) );
  CKND2D0 U3706 ( .A1(n4018), .A2(n4151), .ZN(n3994) );
  OA221D0 U3707 ( .A1(n4152), .A2(n4153), .B1(n4154), .B2(n4155), .C(n4156), 
        .Z(n4018) );
  AOI221D0 U3708 ( .A1(n4157), .A2(n4158), .B1(n4159), .B2(n4160), .C(n3792), 
        .ZN(n4154) );
  IND2D0 U3709 ( .A1(n4161), .B1(n4162), .ZN(n4160) );
  OAI221D0 U3710 ( .A1(n4153), .A2(n4163), .B1(n4164), .B2(n4165), .C(n4166), 
        .ZN(n4158) );
  NR4D0 U3711 ( .A1(n4167), .A2(n4168), .A3(n3807), .A4(n4169), .ZN(n4164) );
  AOI31D0 U3712 ( .A1(n3782), .A2(n3830), .A3(n4170), .B(n4153), .ZN(n4169) );
  NR2D0 U3713 ( .A1(n4171), .A2(n4172), .ZN(n4170) );
  AOI21D0 U3714 ( .A1(n4173), .A2(n4174), .B(n4130), .ZN(n4168) );
  OAI21D0 U3715 ( .A1(n4175), .A2(n4176), .B(n4159), .ZN(n4174) );
  NR3D0 U3716 ( .A1(n3778), .A2(n4177), .A3(n4178), .ZN(n4163) );
  NR3D0 U3717 ( .A1(n4179), .A2(n3773), .A3(n3818), .ZN(n4152) );
  CKND0 U3718 ( .I(n4180), .ZN(n3818) );
  OAI221D0 U3719 ( .A1(n4181), .A2(n4182), .B1(n4183), .B2(n3769), .C(n3814), 
        .ZN(n4046) );
  CKND0 U3720 ( .I(n4143), .ZN(n3814) );
  AOI221D0 U3721 ( .A1(n4184), .A2(n4185), .B1(n3776), .B2(n4186), .C(n4187), 
        .ZN(n4183) );
  OAI221D0 U3722 ( .A1(n4182), .A2(n4188), .B1(n3837), .B2(n4130), .C(n4189), 
        .ZN(n4186) );
  NR4D0 U3723 ( .A1(n4190), .A2(n4135), .A3(n4191), .A4(n4192), .ZN(n4188) );
  ND3D0 U3724 ( .A1(n3600), .A2(n4193), .A3(n3811), .ZN(n4190) );
  IND4D0 U3725 ( .A1(n3799), .B1(n4140), .B2(n4194), .B3(n4195), .ZN(n4185) );
  NR2D0 U3726 ( .A1(n4167), .A2(n3801), .ZN(n4194) );
  ND3D0 U3727 ( .A1(n4196), .A2(n4197), .A3(n4198), .ZN(n3799) );
  NR2D0 U3728 ( .A1(n4142), .A2(n3788), .ZN(n4181) );
  ND3D0 U3729 ( .A1(n4199), .A2(n4200), .A3(n4201), .ZN(n3788) );
  OA221D0 U3730 ( .A1(n4202), .A2(n4203), .B1(n4204), .B2(n3769), .C(n4201), 
        .Z(n3945) );
  CKND0 U3731 ( .I(n4141), .ZN(n4201) );
  OAI21D0 U3732 ( .A1(n4205), .A2(n4206), .B(n4207), .ZN(n4141) );
  CKND2D0 U3733 ( .A1(n4157), .A2(n3771), .ZN(n3769) );
  AOI221D0 U3734 ( .A1(n4208), .A2(n4209), .B1(n3776), .B2(n4210), .C(n4139), 
        .ZN(n4204) );
  CKND2D0 U3735 ( .A1(n4211), .A2(n4196), .ZN(n4139) );
  OAI221D0 U3736 ( .A1(n4203), .A2(n4212), .B1(n4213), .B2(n4130), .C(n4138), 
        .ZN(n4210) );
  AN2D0 U3737 ( .A1(n4214), .A2(n4215), .Z(n4138) );
  AOI21D0 U3738 ( .A1(n4208), .A2(n4216), .B(n4137), .ZN(n4213) );
  CKND2D0 U3739 ( .A1(n4217), .A2(n4218), .ZN(n4137) );
  IND4D0 U3740 ( .A1(n4135), .B1(n3837), .B2(n3838), .B3(n3600), .ZN(n4216) );
  AN2D0 U3741 ( .A1(n4219), .A2(n4220), .Z(n3838) );
  NR2D0 U3742 ( .A1(n3829), .A2(n4134), .ZN(n4212) );
  ND4D0 U3743 ( .A1(n4189), .A2(n4195), .A3(n3323), .A4(n3803), .ZN(n4134) );
  CKND0 U3744 ( .I(n4171), .ZN(n4195) );
  AN2D0 U3745 ( .A1(n3840), .A2(n3834), .Z(n4189) );
  CKND2D0 U3746 ( .A1(n4221), .A2(n4222), .ZN(n3829) );
  CKND0 U3747 ( .I(n4165), .ZN(n3776) );
  ND3D0 U3748 ( .A1(n3822), .A2(n3820), .A3(n4140), .ZN(n4209) );
  INR4D0 U3749 ( .A1(n4223), .B1(n4224), .B2(n3800), .B3(n3292), .ZN(n4140) );
  CKND0 U3750 ( .I(n4129), .ZN(n3820) );
  CKND2D0 U3751 ( .A1(n4197), .A2(n4225), .ZN(n4129) );
  CKND0 U3752 ( .I(n4187), .ZN(n3822) );
  CKND2D0 U3753 ( .A1(n4226), .A2(n4227), .ZN(n4187) );
  NR3D0 U3754 ( .A1(n4143), .A2(n4142), .A3(n4125), .ZN(n4202) );
  OAI21D0 U3755 ( .A1(n4228), .A2(n4200), .B(n4199), .ZN(n4125) );
  ND4D0 U3756 ( .A1(n3287), .A2(n4162), .A3(n4229), .A4(n4230), .ZN(n4142) );
  NR2D0 U3757 ( .A1(n3816), .A2(n3792), .ZN(n4229) );
  NR4D0 U3758 ( .A1(n3789), .A2(n4231), .A3(n3773), .A4(n3817), .ZN(n3287) );
  CKND0 U3759 ( .I(n4232), .ZN(n3817) );
  CKND2D0 U3760 ( .A1(n4233), .A2(n4234), .ZN(n4143) );
  OA221D0 U3761 ( .A1(n4235), .A2(n4236), .B1(n4237), .B2(n4155), .C(n4238), 
        .Z(n4015) );
  AOI221D0 U3762 ( .A1(n4157), .A2(n4239), .B1(n4240), .B2(n4241), .C(n4242), 
        .ZN(n4237) );
  IND2D0 U3763 ( .A1(n3793), .B1(n4243), .ZN(n4241) );
  OAI221D0 U3764 ( .A1(n4236), .A2(n4244), .B1(n4245), .B2(n4165), .C(n4246), 
        .ZN(n4239) );
  CKND0 U3765 ( .I(n3778), .ZN(n4246) );
  AOI221D0 U3766 ( .A1(n3808), .A2(n4247), .B1(n4248), .B2(n4240), .C(n3786), 
        .ZN(n4245) );
  CKND2D0 U3767 ( .A1(n4249), .A2(n3839), .ZN(n4248) );
  OAI221D0 U3768 ( .A1(n4250), .A2(n3810), .B1(n4236), .B2(n4251), .C(n4252), 
        .ZN(n4247) );
  INR4D0 U3769 ( .A1(n3831), .B1(n4253), .B2(n4254), .B3(n4255), .ZN(n4251) );
  IND3D0 U3770 ( .A1(n4256), .B1(n3835), .B2(n3809), .ZN(n4253) );
  NR4D0 U3771 ( .A1(n4257), .A2(n4175), .A3(n3602), .A4(n4192), .ZN(n3809) );
  NR2D0 U3772 ( .A1(n4178), .A2(n4258), .ZN(n4244) );
  NR2D0 U3773 ( .A1(n3789), .A2(n4179), .ZN(n4235) );
  CKND0 U3774 ( .I(n4012), .ZN(n3960) );
  OAI221D0 U3775 ( .A1(n4259), .A2(n4260), .B1(n4261), .B2(n4155), .C(n4180), 
        .ZN(n4012) );
  AOI221D0 U3776 ( .A1(n4157), .A2(n4262), .B1(n4263), .B2(n4264), .C(n3793), 
        .ZN(n4261) );
  CKND2D0 U3777 ( .A1(n4243), .A2(n3775), .ZN(n4264) );
  OAI221D0 U3778 ( .A1(n4260), .A2(n4265), .B1(n4266), .B2(n4165), .C(n4267), 
        .ZN(n4262) );
  INR4D0 U3779 ( .A1(n3804), .B1(n4268), .B2(n3806), .B3(n4269), .ZN(n4266) );
  AOI31D0 U3780 ( .A1(n4270), .A2(n4271), .A3(n4272), .B(n4260), .ZN(n4269) );
  NR3D0 U3781 ( .A1(n3807), .A2(n4273), .A3(n3786), .ZN(n4272) );
  CKND0 U3782 ( .I(n4274), .ZN(n3786) );
  CKND0 U3783 ( .I(n4172), .ZN(n4270) );
  ND3D0 U3784 ( .A1(n4275), .A2(n3831), .A3(n3780), .ZN(n4172) );
  CKND0 U3785 ( .I(n4276), .ZN(n3780) );
  AOI21D0 U3786 ( .A1(n3836), .A2(n4277), .B(n4130), .ZN(n4268) );
  CKND0 U3787 ( .I(n3784), .ZN(n4130) );
  NR2D0 U3788 ( .A1(n3781), .A2(n3810), .ZN(n3784) );
  OAI21D0 U3789 ( .A1(n4257), .A2(n4176), .B(n4263), .ZN(n4277) );
  IND3D0 U3790 ( .A1(n3785), .B1(n3835), .B2(n4278), .ZN(n4176) );
  NR3D0 U3791 ( .A1(n4279), .A2(n3293), .A3(n4224), .ZN(n4265) );
  NR3D0 U3792 ( .A1(n4179), .A2(n3773), .A3(n4280), .ZN(n4259) );
  ND3D0 U3793 ( .A1(n4281), .A2(n4232), .A3(n3289), .ZN(n4179) );
  CKND0 U3794 ( .I(n4282), .ZN(n3289) );
  OAI21D0 U3795 ( .A1(n3894), .A2(n3895), .B(n4283), .ZN(n4020) );
  OAI221D0 U3796 ( .A1(n4284), .A2(n4285), .B1(n4286), .B2(n4155), .C(n4232), 
        .ZN(n3895) );
  CKND2D0 U3797 ( .A1(n4287), .A2(n4281), .ZN(n4232) );
  AOI221D0 U3798 ( .A1(n4157), .A2(n4288), .B1(n4289), .B2(n4290), .C(n3816), 
        .ZN(n4286) );
  ND4D0 U3799 ( .A1(n4162), .A2(n3774), .A3(n4230), .A4(n4291), .ZN(n4290) );
  OAI221D0 U3800 ( .A1(n4285), .A2(n4292), .B1(n4293), .B2(n4165), .C(n4294), 
        .ZN(n4288) );
  CKND0 U3801 ( .I(n4178), .ZN(n4294) );
  CKND2D0 U3802 ( .A1(n3825), .A2(n3824), .ZN(n4178) );
  ND3D0 U3803 ( .A1(n4295), .A2(n4296), .A3(n4297), .ZN(n4165) );
  AOI211D0 U3804 ( .A1(n4298), .A2(n4299), .B(n4300), .C(n4301), .ZN(n4297) );
  OAI22D0 U3805 ( .A1(n4302), .A2(n4208), .B1(n4043), .B2(n4126), .ZN(n4299)
         );
  AOI221D0 U3806 ( .A1(n3808), .A2(n4303), .B1(n4304), .B2(n4289), .C(n4273), 
        .ZN(n4293) );
  CKND0 U3807 ( .I(n3839), .ZN(n4273) );
  CKND2D0 U3808 ( .A1(n4249), .A2(n4274), .ZN(n4304) );
  AN2D0 U3809 ( .A1(n4271), .A2(n3804), .Z(n4249) );
  AN3D0 U3810 ( .A1(n3803), .A2(n4305), .A3(n3782), .Z(n4271) );
  OAI221D0 U3811 ( .A1(n4285), .A2(n4306), .B1(n3835), .B2(n3810), .C(n3831), 
        .ZN(n4303) );
  OAI21D0 U3812 ( .A1(n4307), .A2(n4308), .B(n4309), .ZN(n3810) );
  AOI22D0 U3813 ( .A1(n4123), .A2(n4310), .B1(n4203), .B2(n4097), .ZN(n4307)
         );
  OA21D0 U3814 ( .A1(n4289), .A2(n3937), .B(n4311), .Z(n3835) );
  NR4D0 U3815 ( .A1(n4256), .A2(n4312), .A3(n4276), .A4(n3785), .ZN(n4306) );
  IND4D0 U3816 ( .A1(n4192), .B1(n3837), .B2(n4193), .B3(n4250), .ZN(n3785) );
  NR2D0 U3817 ( .A1(n4313), .A2(n4314), .ZN(n4250) );
  CKND0 U3818 ( .I(n4315), .ZN(n4314) );
  CKND0 U3819 ( .I(n4316), .ZN(n4313) );
  CKND0 U3820 ( .I(n4254), .ZN(n3837) );
  CKND2D0 U3821 ( .A1(n4317), .A2(n3601), .ZN(n4254) );
  CKND2D0 U3822 ( .A1(n3322), .A2(n4252), .ZN(n4276) );
  CKND2D0 U3823 ( .A1(n4173), .A2(n3836), .ZN(n4312) );
  CKND0 U3824 ( .I(n4175), .ZN(n3836) );
  CKND2D0 U3825 ( .A1(n4318), .A2(n4319), .ZN(n4175) );
  CKND0 U3826 ( .I(n4257), .ZN(n4173) );
  CKND2D0 U3827 ( .A1(n4320), .A2(n4321), .ZN(n4257) );
  CKND2D0 U3828 ( .A1(n4322), .A2(n4278), .ZN(n4256) );
  CKND0 U3829 ( .I(n3781), .ZN(n3808) );
  OAI21D0 U3830 ( .A1(n4323), .A2(n4324), .B(n4325), .ZN(n3781) );
  AOI22D0 U3831 ( .A1(n4123), .A2(n4326), .B1(n4203), .B2(n4076), .ZN(n4323)
         );
  NR2D0 U3832 ( .A1(n4258), .A2(n3778), .ZN(n4292) );
  CKND2D0 U3833 ( .A1(n4327), .A2(n4328), .ZN(n3778) );
  IND2D0 U3834 ( .A1(n4177), .B1(n4166), .ZN(n4258) );
  AN2D0 U3835 ( .A1(n3794), .A2(n3795), .Z(n4166) );
  IND4D0 U3836 ( .A1(n3779), .B1(n4267), .B2(n4329), .B3(n4330), .ZN(n4177) );
  NR2D0 U3837 ( .A1(n3800), .A2(n3292), .ZN(n4267) );
  IND2D0 U3838 ( .A1(n4279), .B1(n4331), .ZN(n3779) );
  INR3D0 U3839 ( .A1(n4332), .B1(n4228), .B2(n4206), .ZN(n4157) );
  CKND0 U3840 ( .I(n4205), .ZN(n4228) );
  NR4D0 U3841 ( .A1(n3773), .A2(n4231), .A3(n3789), .A4(n4282), .ZN(n4284) );
  ND3D0 U3842 ( .A1(n4199), .A2(n4207), .A3(n4233), .ZN(n4282) );
  ND4D0 U3843 ( .A1(n4333), .A2(n4182), .A3(n4334), .A4(n4335), .ZN(n4233) );
  NR3D0 U3844 ( .A1(n3372), .A2(n4336), .A3(n4337), .ZN(n4335) );
  ND4D0 U3845 ( .A1(n3771), .A2(n4333), .A3(n4203), .A4(n3946), .ZN(n4207) );
  ND3D0 U3846 ( .A1(n3771), .A2(n4333), .A3(n4338), .ZN(n4199) );
  AOI211D0 U3847 ( .A1(n4203), .A2(n3946), .B(n4126), .C(n3373), .ZN(n4338) );
  CKND0 U3848 ( .I(n4155), .ZN(n3771) );
  OAI211D0 U3849 ( .A1(n4339), .A2(n4340), .B(n4341), .C(n4334), .ZN(n4155) );
  AOI21D0 U3850 ( .A1(n4182), .A2(n4014), .B(n4336), .ZN(n4339) );
  CKND2D0 U3851 ( .A1(n4180), .A2(n4156), .ZN(n3789) );
  CKND0 U3852 ( .I(n4280), .ZN(n4156) );
  NR3D0 U3853 ( .A1(n4287), .A2(n4231), .A3(n4342), .ZN(n4280) );
  CKND2D0 U3854 ( .A1(n4337), .A2(n4334), .ZN(n4180) );
  CKND0 U3855 ( .I(n4238), .ZN(n3773) );
  ND4D0 U3856 ( .A1(n4336), .A2(n4334), .A3(n4333), .A4(n4341), .ZN(n4238) );
  CKND0 U3857 ( .I(n4337), .ZN(n4341) );
  NR3D0 U3858 ( .A1(n4263), .A2(n4011), .A3(n4340), .ZN(n4337) );
  INR3D0 U3859 ( .A1(n4342), .B1(n4231), .B2(n4287), .ZN(n4334) );
  NR3D0 U3860 ( .A1(n3894), .A2(n4289), .A3(n4340), .ZN(n4287) );
  CKND0 U3861 ( .I(n4281), .ZN(n4231) );
  CKND2D0 U3862 ( .A1(n4333), .A2(n3893), .ZN(n4281) );
  ND3D0 U3863 ( .A1(n4153), .A2(n4019), .A3(n4333), .ZN(n4342) );
  CKND0 U3864 ( .I(n4340), .ZN(n4333) );
  CKND2D0 U3865 ( .A1(n3288), .A2(n4343), .ZN(n4340) );
  AN2D0 U3866 ( .A1(n4162), .A2(n4243), .Z(n3288) );
  NR2D0 U3867 ( .A1(n4161), .A2(n3792), .ZN(n4243) );
  CKND0 U3868 ( .I(n4291), .ZN(n3792) );
  CKND2D0 U3869 ( .A1(n4344), .A2(n4345), .ZN(n4291) );
  IND3D0 U3870 ( .A1(n3816), .B1(n4230), .B2(n3774), .ZN(n4161) );
  OA211D0 U3871 ( .A1(n4205), .A2(n4206), .B(n4234), .C(n4200), .Z(n3774) );
  OR2D0 U3872 ( .A1(n4332), .A2(n4206), .Z(n4200) );
  ND3D0 U3873 ( .A1(n4123), .A2(n4028), .A3(n4343), .ZN(n4332) );
  IND3D0 U3874 ( .A1(n4346), .B1(n4347), .B2(n4348), .ZN(n4234) );
  ND3D0 U3875 ( .A1(n4346), .A2(n4348), .A3(n4347), .ZN(n4206) );
  ND3D0 U3876 ( .A1(n4182), .A2(n4029), .A3(n4343), .ZN(n4346) );
  ND3D0 U3877 ( .A1(n4203), .A2(n4034), .A3(n4343), .ZN(n4205) );
  INR2D0 U3878 ( .A1(n4230), .B1(n4349), .ZN(n3816) );
  NR2D0 U3879 ( .A1(n3793), .A2(n4242), .ZN(n4162) );
  CKND0 U3880 ( .I(n3775), .ZN(n4242) );
  IND2D0 U3881 ( .A1(n4348), .B1(n4347), .ZN(n3775) );
  AN3D0 U3882 ( .A1(n4350), .A2(n4351), .A3(n4345), .Z(n4347) );
  ND3D0 U3883 ( .A1(n4236), .A2(n4033), .A3(n4343), .ZN(n4348) );
  INR3D0 U3884 ( .A1(n4345), .B1(n4344), .B2(n4351), .ZN(n3793) );
  ND3D0 U3885 ( .A1(n4260), .A2(n4038), .A3(n4343), .ZN(n4351) );
  CKND0 U3886 ( .I(n4350), .ZN(n4344) );
  ND3D0 U3887 ( .A1(n4153), .A2(n4037), .A3(n4343), .ZN(n4350) );
  AN2D0 U3888 ( .A1(n4349), .A2(n4230), .Z(n4345) );
  CKND2D0 U3889 ( .A1(n4343), .A2(n4035), .ZN(n4230) );
  ND3D0 U3890 ( .A1(n4352), .A2(n4285), .A3(n4343), .ZN(n4349) );
  AN2D0 U3891 ( .A1(n3291), .A2(n4298), .Z(n4343) );
  NR3D0 U3892 ( .A1(n4224), .A2(n3800), .A3(n4279), .ZN(n3291) );
  CKND2D0 U3893 ( .A1(n4198), .A2(n4227), .ZN(n4279) );
  IND3D0 U3894 ( .A1(n4353), .B1(n4354), .B2(n4355), .ZN(n4227) );
  AN2D0 U3895 ( .A1(n4211), .A2(n4225), .Z(n4198) );
  ND3D0 U3896 ( .A1(n4295), .A2(n4298), .A3(n4356), .ZN(n4225) );
  AOI211D0 U3897 ( .A1(n4203), .A2(n4042), .B(n4126), .C(n4043), .ZN(n4356) );
  ND4D0 U3898 ( .A1(n4295), .A2(n4298), .A3(n4203), .A4(n4042), .ZN(n4211) );
  AN3D0 U3899 ( .A1(n4353), .A2(n4355), .A3(n4354), .Z(n4295) );
  ND3D0 U3900 ( .A1(n4182), .A2(n4047), .A3(n4298), .ZN(n4353) );
  CKND0 U3901 ( .I(n3826), .ZN(n3800) );
  IND3D0 U3902 ( .A1(n4357), .B1(n4358), .B2(n4359), .ZN(n3826) );
  ND4D0 U3903 ( .A1(n4329), .A2(n3794), .A3(n4327), .A4(n3825), .ZN(n4224) );
  IND2D0 U3904 ( .A1(n4360), .B1(n4329), .ZN(n3825) );
  IND2D0 U3905 ( .A1(n4355), .B1(n4354), .ZN(n4327) );
  AN3D0 U3906 ( .A1(n4358), .A2(n4357), .A3(n4359), .Z(n4354) );
  ND3D0 U3907 ( .A1(n4260), .A2(n4051), .A3(n4298), .ZN(n4357) );
  ND3D0 U3908 ( .A1(n4236), .A2(n4053), .A3(n4298), .ZN(n4355) );
  IND2D0 U3909 ( .A1(n4358), .B1(n4359), .ZN(n3794) );
  AN2D0 U3910 ( .A1(n4360), .A2(n4329), .Z(n4359) );
  ND3D0 U3911 ( .A1(n4361), .A2(n4285), .A3(n4298), .ZN(n4360) );
  ND3D0 U3912 ( .A1(n4153), .A2(n4052), .A3(n4298), .ZN(n4358) );
  CKND2D0 U3913 ( .A1(n4298), .A2(n4049), .ZN(n4329) );
  INR3D0 U3914 ( .A1(n4362), .B1(n3293), .B2(n3292), .ZN(n4298) );
  CKND0 U3915 ( .I(n3796), .ZN(n3292) );
  IND3D0 U3916 ( .A1(n4363), .B1(n4364), .B2(n4365), .ZN(n3796) );
  CKND2D0 U3917 ( .A1(n4223), .A2(n4331), .ZN(n3293) );
  AN3D0 U3918 ( .A1(n4226), .A2(n4197), .A3(n4196), .Z(n4331) );
  CKND2D0 U3919 ( .A1(n4300), .A2(n4296), .ZN(n4196) );
  CKND0 U3920 ( .I(n4366), .ZN(n4300) );
  ND3D0 U3921 ( .A1(n4301), .A2(n4366), .A3(n4296), .ZN(n4197) );
  AN3D0 U3922 ( .A1(n4367), .A2(n4368), .A3(n4369), .Z(n4296) );
  ND3D0 U3923 ( .A1(n4203), .A2(n4062), .A3(n4362), .ZN(n4366) );
  AN3D0 U3924 ( .A1(n4123), .A2(n4060), .A3(n4362), .Z(n4301) );
  IND3D0 U3925 ( .A1(n4368), .B1(n4369), .B2(n4367), .ZN(n4226) );
  ND3D0 U3926 ( .A1(n4182), .A2(n4065), .A3(n4362), .ZN(n4368) );
  AN4D0 U3927 ( .A1(n4330), .A2(n3795), .A3(n4328), .A4(n3824), .Z(n4223) );
  IND2D0 U3928 ( .A1(n4370), .B1(n4330), .ZN(n3824) );
  IND2D0 U3929 ( .A1(n4367), .B1(n4369), .ZN(n4328) );
  AN3D0 U3930 ( .A1(n4364), .A2(n4363), .A3(n4365), .Z(n4369) );
  ND3D0 U3931 ( .A1(n4260), .A2(n4070), .A3(n4362), .ZN(n4363) );
  ND3D0 U3932 ( .A1(n4236), .A2(n4066), .A3(n4362), .ZN(n4367) );
  IND2D0 U3933 ( .A1(n4364), .B1(n4365), .ZN(n3795) );
  AN2D0 U3934 ( .A1(n4370), .A2(n4330), .Z(n4365) );
  ND3D0 U3935 ( .A1(n4371), .A2(n4285), .A3(n4362), .ZN(n4370) );
  ND3D0 U3936 ( .A1(n4153), .A2(n4069), .A3(n4362), .ZN(n4364) );
  CKND2D0 U3937 ( .A1(n4362), .A2(n4067), .ZN(n4330) );
  INR2D0 U3938 ( .A1(n3603), .B1(n4324), .ZN(n4362) );
  INR3D0 U3939 ( .A1(n3782), .B1(n4167), .B2(n4171), .ZN(n3603) );
  ND4D0 U3940 ( .A1(n3804), .A2(n4305), .A3(n4274), .A4(n3839), .ZN(n4171) );
  CKND2D0 U3941 ( .A1(n4372), .A2(n4305), .ZN(n3839) );
  CKND2D0 U3942 ( .A1(n4373), .A2(n4374), .ZN(n4274) );
  ND3D0 U3943 ( .A1(n4375), .A2(n4376), .A3(n4377), .ZN(n3804) );
  CKND0 U3944 ( .I(n3803), .ZN(n4167) );
  CKND2D0 U3945 ( .A1(n4378), .A2(n4375), .ZN(n3803) );
  INR2D0 U3946 ( .A1(n3840), .B1(n3801), .ZN(n3782) );
  CKND2D0 U3947 ( .A1(n4215), .A2(n4222), .ZN(n3801) );
  ND3D0 U3948 ( .A1(n4325), .A2(n4379), .A3(n4380), .ZN(n4222) );
  AOI211D0 U3949 ( .A1(n4203), .A2(n4076), .B(n4126), .C(n4077), .ZN(n4380) );
  ND4D0 U3950 ( .A1(n4325), .A2(n4379), .A3(n4203), .A4(n4076), .ZN(n4215) );
  INR3D0 U3951 ( .A1(n4373), .B1(n4381), .B2(n4374), .ZN(n4325) );
  CKND0 U3952 ( .I(n4382), .ZN(n4374) );
  ND3D0 U3953 ( .A1(n4373), .A2(n4382), .A3(n4381), .ZN(n3840) );
  NR3D0 U3954 ( .A1(n4184), .A2(n4074), .A3(n4324), .ZN(n4381) );
  ND3D0 U3955 ( .A1(n4236), .A2(n4083), .A3(n4379), .ZN(n4382) );
  INR3D0 U3956 ( .A1(n4375), .B1(n4377), .B2(n4378), .ZN(n4373) );
  CKND0 U3957 ( .I(n4376), .ZN(n4378) );
  ND3D0 U3958 ( .A1(n4153), .A2(n4082), .A3(n4379), .ZN(n4376) );
  NR3D0 U3959 ( .A1(n4263), .A2(n4004), .A3(n4324), .ZN(n4377) );
  INR2D0 U3960 ( .A1(n4305), .B1(n4372), .ZN(n4375) );
  NR3D0 U3961 ( .A1(n4080), .A2(n4289), .A3(n4324), .ZN(n4372) );
  CKND2D0 U3962 ( .A1(n4379), .A2(n4079), .ZN(n4305) );
  CKND0 U3963 ( .I(n4324), .ZN(n4379) );
  ND3D0 U3964 ( .A1(n4383), .A2(n3323), .A3(n3322), .ZN(n4324) );
  CKND0 U3965 ( .I(n4255), .ZN(n3322) );
  CKND2D0 U3966 ( .A1(n3811), .A2(n3834), .ZN(n4255) );
  IND3D0 U3967 ( .A1(n4384), .B1(n4385), .B2(n4386), .ZN(n3834) );
  AN2D0 U3968 ( .A1(n4214), .A2(n4221), .Z(n3811) );
  ND3D0 U3969 ( .A1(n4309), .A2(n4383), .A3(n4387), .ZN(n4221) );
  AOI211D0 U3970 ( .A1(n4203), .A2(n4097), .B(n4126), .C(n4092), .ZN(n4387) );
  ND4D0 U3971 ( .A1(n4309), .A2(n4383), .A3(n4203), .A4(n4097), .ZN(n4214) );
  AN3D0 U3972 ( .A1(n4384), .A2(n4386), .A3(n4385), .Z(n4309) );
  ND3D0 U3973 ( .A1(n4182), .A2(n4087), .A3(n4383), .ZN(n4384) );
  CKND0 U3974 ( .I(n4191), .ZN(n3323) );
  ND3D0 U3975 ( .A1(n4252), .A2(n3831), .A3(n4322), .ZN(n4191) );
  INR3D0 U3976 ( .A1(n4275), .B1(n3806), .B2(n3807), .ZN(n4322) );
  INR2D0 U3977 ( .A1(n4388), .B1(n4389), .ZN(n3807) );
  CKND0 U3978 ( .I(n3830), .ZN(n3806) );
  IND3D0 U3979 ( .A1(n4390), .B1(n4388), .B2(n4389), .ZN(n3830) );
  CKND2D0 U3980 ( .A1(n4391), .A2(n4275), .ZN(n3831) );
  IND2D0 U3981 ( .A1(n4386), .B1(n4385), .ZN(n4252) );
  AN3D0 U3982 ( .A1(n4389), .A2(n4390), .A3(n4388), .Z(n4385) );
  INR2D0 U3983 ( .A1(n4275), .B1(n4391), .ZN(n4388) );
  NR3D0 U3984 ( .A1(n4099), .A2(n4289), .A3(n4308), .ZN(n4391) );
  CKND2D0 U3985 ( .A1(n4383), .A2(n4098), .ZN(n4275) );
  ND3D0 U3986 ( .A1(n4260), .A2(n4101), .A3(n4383), .ZN(n4390) );
  ND3D0 U3987 ( .A1(n4153), .A2(n4100), .A3(n4383), .ZN(n4389) );
  ND3D0 U3988 ( .A1(n4236), .A2(n4096), .A3(n4383), .ZN(n4386) );
  CKND0 U3989 ( .I(n4308), .ZN(n4383) );
  ND4D0 U3990 ( .A1(n3600), .A2(n4193), .A3(n4392), .A4(n3601), .ZN(n4308) );
  ND3D0 U3991 ( .A1(n4393), .A2(n4392), .A3(n4394), .ZN(n3601) );
  AOI211D0 U3992 ( .A1(n4236), .A2(n4115), .B(n4184), .C(n4114), .ZN(n4394) );
  CKND0 U3993 ( .I(n3602), .ZN(n4193) );
  CKND2D0 U3994 ( .A1(n4218), .A2(n4220), .ZN(n3602) );
  ND3D0 U3995 ( .A1(n4395), .A2(n4392), .A3(n4396), .ZN(n4220) );
  AOI211D0 U3996 ( .A1(n4203), .A2(n4106), .B(n4126), .C(n4107), .ZN(n4396) );
  ND4D0 U3997 ( .A1(n4395), .A2(n4392), .A3(n4203), .A4(n4106), .ZN(n4218) );
  OA221D0 U3998 ( .A1(n4397), .A2(n4240), .B1(n4114), .B2(n4184), .C(n4393), 
        .Z(n4395) );
  CKND0 U3999 ( .I(n4136), .ZN(n3600) );
  ND4D0 U4000 ( .A1(n4311), .A2(n4278), .A3(n4315), .A4(n4398), .ZN(n4136) );
  AN2D0 U4001 ( .A1(n4319), .A2(n4320), .Z(n4398) );
  IND2D0 U4002 ( .A1(n4399), .B1(n4400), .ZN(n4320) );
  IND3D0 U4003 ( .A1(n4401), .B1(n4400), .B2(n4399), .ZN(n4319) );
  ND4D0 U4004 ( .A1(n4393), .A2(n4392), .A3(n4236), .A4(n4115), .ZN(n4315) );
  CKND0 U4005 ( .I(n4240), .ZN(n4236) );
  AN3D0 U4006 ( .A1(n4399), .A2(n4401), .A3(n4400), .Z(n4393) );
  AN2D0 U4007 ( .A1(n4402), .A2(n4278), .Z(n4400) );
  ND3D0 U4008 ( .A1(n4260), .A2(n4104), .A3(n4392), .ZN(n4401) );
  CKND0 U4009 ( .I(n4263), .ZN(n4260) );
  ND3D0 U4010 ( .A1(n4153), .A2(n4113), .A3(n4392), .ZN(n4399) );
  IND2D0 U4011 ( .A1(n4402), .B1(n4278), .ZN(n4311) );
  CKND2D0 U4012 ( .A1(n4392), .A2(n4112), .ZN(n4278) );
  ND3D0 U4013 ( .A1(n4111), .A2(n4285), .A3(n4392), .ZN(n4402) );
  INR3D0 U4014 ( .A1(n4317), .B1(n4192), .B2(n4135), .ZN(n4392) );
  ND4D0 U4015 ( .A1(n4318), .A2(n4150), .A3(n4316), .A4(n4403), .ZN(n4135) );
  OA21D0 U4016 ( .A1(n3937), .A2(n4289), .B(n4321), .Z(n4403) );
  CKND2D0 U4017 ( .A1(n4404), .A2(n4405), .ZN(n4321) );
  IND4D0 U4018 ( .A1(n4406), .B1(n4407), .B2(n4405), .B3(n4408), .ZN(n4316) );
  ND3D0 U4019 ( .A1(n4405), .A2(n4408), .A3(n4406), .ZN(n4318) );
  CKND2D0 U4020 ( .A1(n4219), .A2(n4217), .ZN(n4192) );
  ND3D0 U4021 ( .A1(n4409), .A2(n4121), .A3(n4203), .ZN(n4217) );
  ND4D0 U4022 ( .A1(n4123), .A2(n4409), .A3(n4119), .A4(n4410), .ZN(n4219) );
  CKND2D0 U4023 ( .A1(n4203), .A2(n4121), .ZN(n4410) );
  CKND0 U4024 ( .I(n4208), .ZN(n4203) );
  OAI221D0 U4025 ( .A1(n4411), .A2(n4412), .B1(n4413), .B2(n3720), .C(n4414), 
        .ZN(n4208) );
  CKND0 U4026 ( .I(n4415), .ZN(n4414) );
  AOI221D0 U4027 ( .A1(n4416), .A2(n4417), .B1(n4418), .B2(n4419), .C(n4420), 
        .ZN(n4413) );
  OAI21D0 U4028 ( .A1(n4421), .A2(n4411), .B(n4422), .ZN(n4419) );
  NR4D0 U4029 ( .A1(n4423), .A2(n3347), .A3(n3754), .A4(n3751), .ZN(n4421) );
  IND2D0 U4030 ( .A1(n3745), .B1(n4424), .ZN(n4416) );
  NR2D0 U4031 ( .A1(n4425), .A2(n4426), .ZN(n4412) );
  OA21D0 U4032 ( .A1(n4146), .A2(n4184), .B(n4427), .Z(n4409) );
  CKND0 U4033 ( .I(n4126), .ZN(n4123) );
  OAI221D0 U4034 ( .A1(n4428), .A2(n4429), .B1(n4430), .B2(n3720), .C(n4431), 
        .ZN(n4126) );
  CKND0 U4035 ( .I(n4425), .ZN(n4431) );
  OAI21D0 U4036 ( .A1(n3737), .A2(n3722), .B(n4432), .ZN(n4425) );
  AN2D0 U4037 ( .A1(n4433), .A2(n4434), .Z(n3737) );
  AOI221D0 U4038 ( .A1(n4418), .A2(n3751), .B1(n4435), .B2(n4436), .C(n3745), 
        .ZN(n4430) );
  CKND2D0 U4039 ( .A1(n4437), .A2(n4438), .ZN(n3745) );
  IND4D0 U4040 ( .A1(n4420), .B1(n4422), .B2(n4424), .B3(n4439), .ZN(n4435) );
  NR3D0 U4041 ( .A1(n3754), .A2(n4423), .A3(n3347), .ZN(n4439) );
  INR4D0 U4042 ( .A1(n3314), .B1(n4440), .B2(n4441), .B3(n4442), .ZN(n4424) );
  AN2D0 U4043 ( .A1(n4443), .A2(n4444), .Z(n4422) );
  CKND2D0 U4044 ( .A1(n4445), .A2(n4446), .ZN(n4420) );
  CKND2D0 U4045 ( .A1(n4447), .A2(n4448), .ZN(n3751) );
  NR2D0 U4046 ( .A1(n4426), .A2(n4415), .ZN(n4429) );
  CKND2D0 U4047 ( .A1(n4449), .A2(n4450), .ZN(n4415) );
  AO21D0 U4048 ( .A1(n4451), .A2(n4452), .B(n3722), .Z(n4450) );
  OAI211D0 U4049 ( .A1(n4453), .A2(n3722), .B(n4454), .C(n4455), .ZN(n4426) );
  ND3D0 U4050 ( .A1(n4182), .A2(n4144), .A3(n4427), .ZN(n4317) );
  INR4D0 U4051 ( .A1(n4405), .B1(n4406), .B2(n4407), .B3(n4404), .ZN(n4427) );
  CKND0 U4052 ( .I(n4408), .ZN(n4404) );
  CKND2D0 U4053 ( .A1(n4153), .A2(n4151), .ZN(n4408) );
  NR2D0 U4054 ( .A1(n4240), .A2(n4456), .ZN(n4407) );
  NR2D0 U4055 ( .A1(n4263), .A2(n4457), .ZN(n4406) );
  OAI221D0 U4056 ( .A1(n4458), .A2(n4459), .B1(n4460), .B2(n3722), .C(n4461), 
        .ZN(n4263) );
  AOI221D0 U4057 ( .A1(n4462), .A2(n4463), .B1(n3699), .B2(n4464), .C(n4465), 
        .ZN(n4460) );
  ND4D0 U4058 ( .A1(n4466), .A2(n3709), .A3(n4467), .A4(n3707), .ZN(n4464) );
  OAI21D0 U4059 ( .A1(n4468), .A2(n3752), .B(n4418), .ZN(n4467) );
  AOI21D0 U4060 ( .A1(n4469), .A2(n4470), .B(n4458), .ZN(n4468) );
  OAI31D0 U4061 ( .A1(n4471), .A2(n4472), .A3(n4473), .B(n4463), .ZN(n4466) );
  ND3D0 U4062 ( .A1(n4474), .A2(n3756), .A3(n3710), .ZN(n4471) );
  ND3D0 U4063 ( .A1(n4475), .A2(n4476), .A3(n4477), .ZN(n4462) );
  NR2D0 U4064 ( .A1(n4478), .A2(n3715), .ZN(n4459) );
  CKND2D0 U4065 ( .A1(n4479), .A2(n4285), .ZN(n4405) );
  CKND0 U4066 ( .I(n4184), .ZN(n4182) );
  OAI211D0 U4067 ( .A1(n4480), .A2(n4481), .B(n4455), .C(n4482), .ZN(n4184) );
  AOI21D0 U4068 ( .A1(n4483), .A2(n4484), .B(n4442), .ZN(n4482) );
  OAI21D0 U4069 ( .A1(n4485), .A2(n3713), .B(n3746), .ZN(n4484) );
  OA211D0 U4070 ( .A1(n3739), .A2(n3722), .B(n3729), .C(n3732), .Z(n4455) );
  AN2D0 U4071 ( .A1(n4486), .A2(n4487), .Z(n3739) );
  NR4D0 U4072 ( .A1(n4488), .A2(n4489), .A3(n3704), .A4(n4440), .ZN(n4481) );
  OAI21D0 U4073 ( .A1(n4490), .A2(n3718), .B(n3706), .ZN(n4489) );
  CKND0 U4074 ( .I(n4483), .ZN(n3718) );
  NR2D0 U4075 ( .A1(n3720), .A2(n3711), .ZN(n4483) );
  CKND2D0 U4076 ( .A1(n3691), .A2(n3699), .ZN(n3720) );
  CKND0 U4077 ( .I(n3722), .ZN(n3691) );
  NR4D0 U4078 ( .A1(n4491), .A2(n4492), .A3(n3347), .A4(n4493), .ZN(n4490) );
  ND3D0 U4079 ( .A1(n4494), .A2(n4495), .A3(n3349), .ZN(n4491) );
  IIND4D0 U4080 ( .A1(n3693), .A2(n3701), .B1(n4453), .B2(n4454), .ZN(n4488)
         );
  AN2D0 U4081 ( .A1(n3269), .A2(n4496), .Z(n4454) );
  AN4D0 U4082 ( .A1(n3734), .A2(n4497), .A3(n3687), .A4(n4498), .Z(n3269) );
  NR2D0 U4083 ( .A1(n4499), .A2(n3694), .ZN(n4498) );
  AN4D0 U4084 ( .A1(n4500), .A2(n4501), .A3(n4502), .A4(n4503), .Z(n4453) );
  ND3D0 U4085 ( .A1(n4451), .A2(n4433), .A3(n4504), .ZN(n3701) );
  CKND2D0 U4086 ( .A1(n4432), .A2(n4449), .ZN(n3693) );
  OA21D0 U4087 ( .A1(n4505), .A2(n4506), .B(n4507), .Z(n4449) );
  CKND0 U4088 ( .I(n3736), .ZN(n4432) );
  CKND2D0 U4089 ( .A1(n4508), .A2(n4509), .ZN(n3736) );
  CKND0 U4090 ( .I(n4289), .ZN(n4285) );
  OAI221D0 U4091 ( .A1(n4510), .A2(n4511), .B1(n4512), .B2(n3722), .C(n4513), 
        .ZN(n4289) );
  AOI221D0 U4092 ( .A1(n4514), .A2(n4515), .B1(n3699), .B2(n4516), .C(n4517), 
        .ZN(n4512) );
  OAI221D0 U4093 ( .A1(n4510), .A2(n4518), .B1(n4519), .B2(n3711), .C(n3756), 
        .ZN(n4516) );
  AOI221D0 U4094 ( .A1(n3725), .A2(n3753), .B1(n4520), .B2(n4515), .C(n4521), 
        .ZN(n4519) );
  ND4D0 U4095 ( .A1(n4522), .A2(n4469), .A3(n4523), .A4(n4524), .ZN(n4520) );
  NR2D0 U4096 ( .A1(n4525), .A2(n3726), .ZN(n4523) );
  NR2D0 U4097 ( .A1(n3723), .A2(n4526), .ZN(n4518) );
  CKND0 U4098 ( .I(n4474), .ZN(n3723) );
  CKND2D0 U4099 ( .A1(n4477), .A2(n4527), .ZN(n4514) );
  CKND0 U4100 ( .I(n4528), .ZN(n4477) );
  INR3D0 U4101 ( .A1(n4529), .B1(n4530), .B2(n4531), .ZN(n4511) );
  CKND0 U4102 ( .I(n4159), .ZN(n4153) );
  OAI221D0 U4103 ( .A1(n4532), .A2(n4533), .B1(n4534), .B2(n3722), .C(n4535), 
        .ZN(n4159) );
  CKND0 U4104 ( .I(n4530), .ZN(n4535) );
  AOI221D0 U4105 ( .A1(n4536), .A2(n4537), .B1(n3699), .B2(n4538), .C(n4528), 
        .ZN(n4534) );
  CKND2D0 U4106 ( .A1(n3695), .A2(n3696), .ZN(n4528) );
  OAI211D0 U4107 ( .A1(n4532), .A2(n4539), .B(n3710), .C(n4540), .ZN(n4538) );
  AOI21D0 U4108 ( .A1(n4418), .A2(n4541), .B(n4441), .ZN(n4540) );
  CKND2D0 U4109 ( .A1(n4469), .A2(n4542), .ZN(n4541) );
  AO21D0 U4110 ( .A1(n4470), .A2(n4524), .B(n4532), .Z(n4542) );
  INR3D0 U4111 ( .A1(n4543), .B1(n3753), .B2(n3726), .ZN(n4470) );
  ND4D0 U4112 ( .A1(n4485), .A2(n3349), .A3(n4544), .A4(n4495), .ZN(n3726) );
  AN2D0 U4113 ( .A1(n4545), .A2(n4546), .Z(n4544) );
  CKND0 U4114 ( .I(n3754), .ZN(n4485) );
  NR2D0 U4115 ( .A1(n3711), .A2(n3713), .ZN(n4418) );
  NR4D0 U4116 ( .A1(n3750), .A2(n3724), .A3(n4440), .A4(n4472), .ZN(n4539) );
  IND3D0 U4117 ( .A1(n3727), .B1(n4547), .B2(n3747), .ZN(n4472) );
  ND3D0 U4118 ( .A1(n3746), .A2(n4548), .A3(n3313), .ZN(n3727) );
  CKND0 U4119 ( .I(n3709), .ZN(n3750) );
  CKND2D0 U4120 ( .A1(n4475), .A2(n4527), .ZN(n4536) );
  INR2D0 U4121 ( .A1(n4476), .B1(n4465), .ZN(n4527) );
  CKND2D0 U4122 ( .A1(n3703), .A2(n3697), .ZN(n4465) );
  AN3D0 U4123 ( .A1(n4549), .A2(n4550), .A3(n3721), .Z(n4476) );
  AN3D0 U4124 ( .A1(n4551), .A2(n4552), .A3(n4553), .Z(n3721) );
  CKND0 U4125 ( .I(n4554), .ZN(n4551) );
  CKND0 U4126 ( .I(n4517), .ZN(n4475) );
  CKND2D0 U4127 ( .A1(n3742), .A2(n3741), .ZN(n4517) );
  NR2D0 U4128 ( .A1(n4555), .A2(n4531), .ZN(n4533) );
  ND3D0 U4129 ( .A1(n3728), .A2(n4497), .A3(n4556), .ZN(n4531) );
  INR2D0 U4130 ( .A1(n4016), .B1(n4240), .ZN(n4336) );
  OAI221D0 U4131 ( .A1(n4557), .A2(n4558), .B1(n4559), .B2(n3722), .C(n4560), 
        .ZN(n4240) );
  CKND0 U4132 ( .I(n3715), .ZN(n4560) );
  CKND2D0 U4133 ( .A1(n4497), .A2(n4561), .ZN(n3715) );
  ND4D0 U4134 ( .A1(n4562), .A2(n4563), .A3(n4564), .A4(n4565), .ZN(n4497) );
  ND4D0 U4135 ( .A1(n4566), .A2(n4567), .A3(n4568), .A4(n4506), .ZN(n3722) );
  AOI221D0 U4136 ( .A1(n4569), .A2(n4570), .B1(n3699), .B2(n4571), .C(n4554), 
        .ZN(n4559) );
  CKND2D0 U4137 ( .A1(n4502), .A2(n4503), .ZN(n4554) );
  OAI221D0 U4138 ( .A1(n4557), .A2(n4572), .B1(n4573), .B2(n3711), .C(n4474), 
        .ZN(n4571) );
  OAI21D0 U4139 ( .A1(n4574), .A2(n4575), .B(n4576), .ZN(n3711) );
  AOI22D0 U4140 ( .A1(n4428), .A2(n4326), .B1(n4411), .B2(n4076), .ZN(n4574)
         );
  AOI221D0 U4141 ( .A1(n4577), .A2(n4570), .B1(n3725), .B2(n4578), .C(n4525), 
        .ZN(n4573) );
  CKND0 U4142 ( .I(n4548), .ZN(n4525) );
  CKND2D0 U4143 ( .A1(n4545), .A2(n4546), .ZN(n4578) );
  CKND0 U4144 ( .I(n3713), .ZN(n3725) );
  OAI21D0 U4145 ( .A1(n4579), .A2(n4580), .B(n4581), .ZN(n3713) );
  AOI22D0 U4146 ( .A1(n4428), .A2(n4310), .B1(n4411), .B2(n4097), .ZN(n4579)
         );
  IND4D0 U4147 ( .A1(n3753), .B1(n3712), .B2(n4522), .B3(n4582), .ZN(n4577) );
  NR2D0 U4148 ( .A1(n4521), .A2(n3754), .ZN(n4582) );
  CKND2D0 U4149 ( .A1(n4583), .A2(n3348), .ZN(n3754) );
  CKND0 U4150 ( .I(n3747), .ZN(n4521) );
  AN4D0 U4151 ( .A1(n3313), .A2(n4584), .A3(n3746), .A4(n4543), .Z(n4522) );
  AN4D0 U4152 ( .A1(n4469), .A2(n4524), .A3(n3349), .A4(n4495), .Z(n3712) );
  CKND0 U4153 ( .I(n3752), .ZN(n4524) );
  CKND2D0 U4154 ( .A1(n4585), .A2(n4586), .ZN(n3752) );
  AN2D0 U4155 ( .A1(n4587), .A2(n4588), .Z(n4469) );
  OAI21D0 U4156 ( .A1(n4515), .A2(n3937), .B(n4589), .ZN(n3753) );
  INR2D0 U4157 ( .A1(n3756), .B1(n4526), .ZN(n4572) );
  IND2D0 U4158 ( .A1(n4473), .B1(n3707), .ZN(n4526) );
  ND3D0 U4159 ( .A1(n3706), .A2(n4590), .A3(n4591), .ZN(n4473) );
  AN3D0 U4160 ( .A1(n4592), .A2(n4593), .A3(n4594), .Z(n3699) );
  AOI211D0 U4161 ( .A1(n4595), .A2(n4596), .B(n4597), .C(n4598), .ZN(n4594) );
  OAI22D0 U4162 ( .A1(n4302), .A2(n4417), .B1(n4043), .B2(n4436), .ZN(n4596)
         );
  IND3D0 U4163 ( .A1(n3273), .B1(n4500), .B2(n4552), .ZN(n4569) );
  INR2D0 U4164 ( .A1(n4461), .B1(n4478), .ZN(n4558) );
  OR2D0 U4165 ( .A1(n4555), .A2(n4530), .Z(n4478) );
  CKND2D0 U4166 ( .A1(n3687), .A2(n3688), .ZN(n4530) );
  IND3D0 U4167 ( .A1(n4599), .B1(n4600), .B2(n4601), .ZN(n3687) );
  CKND2D0 U4168 ( .A1(n4513), .A2(n4529), .ZN(n4555) );
  INR3D0 U4169 ( .A1(n4602), .B1(n4499), .B2(n3714), .ZN(n4529) );
  CKND2D0 U4170 ( .A1(n3267), .A2(n4603), .ZN(n3714) );
  AN3D0 U4171 ( .A1(n3729), .A2(n4507), .A3(n4509), .Z(n3267) );
  ND3D0 U4172 ( .A1(n4566), .A2(n4564), .A3(n4604), .ZN(n4509) );
  AOI211D0 U4173 ( .A1(n4411), .A2(n3946), .B(n4436), .C(n3373), .ZN(n4604) );
  ND4D0 U4174 ( .A1(n4566), .A2(n4564), .A3(n4411), .A4(n3946), .ZN(n4507) );
  OA211D0 U4175 ( .A1(n4605), .A2(n4606), .B(n4565), .C(n4563), .Z(n4566) );
  CKND0 U4176 ( .I(n4607), .ZN(n4565) );
  AOI21D0 U4177 ( .A1(n4480), .A2(n4014), .B(n4562), .ZN(n4605) );
  ND4D0 U4178 ( .A1(n4564), .A2(n4480), .A3(n4563), .A4(n4608), .ZN(n3729) );
  NR3D0 U4179 ( .A1(n3372), .A2(n4562), .A3(n4607), .ZN(n4608) );
  INR2D0 U4180 ( .A1(n4016), .B1(n4570), .ZN(n4562) );
  AN2D0 U4181 ( .A1(n3734), .A2(n3733), .Z(n4513) );
  OR2D0 U4182 ( .A1(n4600), .A2(n4499), .Z(n3734) );
  CKND0 U4183 ( .I(n4601), .ZN(n4499) );
  INR2D0 U4184 ( .A1(n3689), .B1(n3694), .ZN(n4461) );
  CKND0 U4185 ( .I(n3728), .ZN(n3694) );
  CKND2D0 U4186 ( .A1(n4607), .A2(n4563), .ZN(n3728) );
  AN3D0 U4187 ( .A1(n4599), .A2(n4601), .A3(n4600), .Z(n4563) );
  IND3D0 U4188 ( .A1(n3894), .B1(n4510), .B2(n4564), .ZN(n4600) );
  CKND2D0 U4189 ( .A1(n4564), .A2(n3893), .ZN(n4601) );
  ND3D0 U4190 ( .A1(n4532), .A2(n4019), .A3(n4564), .ZN(n4599) );
  CKND0 U4191 ( .I(n4606), .ZN(n4564) );
  NR3D0 U4192 ( .A1(n4463), .A2(n4011), .A3(n4606), .ZN(n4607) );
  CKND2D0 U4193 ( .A1(n3268), .A2(n4609), .ZN(n4606) );
  AN2D0 U4194 ( .A1(n4496), .A2(n4603), .Z(n3268) );
  OA211D0 U4195 ( .A1(n4505), .A2(n4506), .B(n3732), .C(n4508), .Z(n4603) );
  IND3D0 U4196 ( .A1(n4568), .B1(n4506), .B2(n4567), .ZN(n4508) );
  CKND0 U4197 ( .I(n4505), .ZN(n4567) );
  ND3D0 U4198 ( .A1(n4428), .A2(n4028), .A3(n4609), .ZN(n4568) );
  IND3D0 U4199 ( .A1(n4610), .B1(n4611), .B2(n4612), .ZN(n3732) );
  ND3D0 U4200 ( .A1(n4411), .A2(n4034), .A3(n4609), .ZN(n4506) );
  ND3D0 U4201 ( .A1(n4610), .A2(n4612), .A3(n4611), .ZN(n4505) );
  ND3D0 U4202 ( .A1(n4480), .A2(n4029), .A3(n4609), .ZN(n4610) );
  AN4D0 U4203 ( .A1(n4556), .A2(n4602), .A3(n3688), .A4(n3733), .Z(n4496) );
  IND2D0 U4204 ( .A1(n4613), .B1(n4602), .ZN(n3733) );
  IND2D0 U4205 ( .A1(n4614), .B1(n4615), .ZN(n3688) );
  AN2D0 U4206 ( .A1(n4561), .A2(n3689), .Z(n4556) );
  IND2D0 U4207 ( .A1(n4612), .B1(n4611), .ZN(n4561) );
  AN3D0 U4208 ( .A1(n4614), .A2(n4616), .A3(n4615), .Z(n4611) );
  ND3D0 U4209 ( .A1(n4557), .A2(n4033), .A3(n4609), .ZN(n4612) );
  IND3D0 U4210 ( .A1(n4616), .B1(n4615), .B2(n4614), .ZN(n3689) );
  ND3D0 U4211 ( .A1(n4532), .A2(n4037), .A3(n4609), .ZN(n4614) );
  AN2D0 U4212 ( .A1(n4613), .A2(n4602), .Z(n4615) );
  CKND2D0 U4213 ( .A1(n4609), .A2(n4035), .ZN(n4602) );
  ND3D0 U4214 ( .A1(n4352), .A2(n4510), .A3(n4609), .ZN(n4613) );
  ND3D0 U4215 ( .A1(n4458), .A2(n4038), .A3(n4609), .ZN(n4616) );
  INR2D0 U4216 ( .A1(n4595), .B1(n3271), .ZN(n4609) );
  ND3D0 U4217 ( .A1(n4500), .A2(n4502), .A3(n4552), .ZN(n3271) );
  AN2D0 U4218 ( .A1(n4504), .A2(n4487), .Z(n4552) );
  IND3D0 U4219 ( .A1(n4617), .B1(n4618), .B2(n4619), .ZN(n4487) );
  AN2D0 U4220 ( .A1(n4452), .A2(n4434), .Z(n4504) );
  ND3D0 U4221 ( .A1(n4592), .A2(n4595), .A3(n4620), .ZN(n4434) );
  AOI211D0 U4222 ( .A1(n4411), .A2(n4042), .B(n4436), .C(n4043), .ZN(n4620) );
  ND4D0 U4223 ( .A1(n4592), .A2(n4595), .A3(n4411), .A4(n4042), .ZN(n4452) );
  AN3D0 U4224 ( .A1(n4617), .A2(n4619), .A3(n4618), .Z(n4592) );
  ND3D0 U4225 ( .A1(n4480), .A2(n4047), .A3(n4595), .ZN(n4617) );
  IND2D0 U4226 ( .A1(n4619), .B1(n4618), .ZN(n4502) );
  AN3D0 U4227 ( .A1(n4621), .A2(n4622), .A3(n4623), .Z(n4618) );
  ND3D0 U4228 ( .A1(n4557), .A2(n4053), .A3(n4595), .ZN(n4619) );
  AN4D0 U4229 ( .A1(n3703), .A2(n4549), .A3(n3695), .A4(n3742), .Z(n4500) );
  IND2D0 U4230 ( .A1(n4624), .B1(n4549), .ZN(n3742) );
  IND2D0 U4231 ( .A1(n4621), .B1(n4623), .ZN(n3695) );
  IND3D0 U4232 ( .A1(n4622), .B1(n4623), .B2(n4621), .ZN(n3703) );
  ND3D0 U4233 ( .A1(n4532), .A2(n4052), .A3(n4595), .ZN(n4621) );
  AN2D0 U4234 ( .A1(n4624), .A2(n4549), .Z(n4623) );
  CKND2D0 U4235 ( .A1(n4595), .A2(n4049), .ZN(n4549) );
  ND3D0 U4236 ( .A1(n4361), .A2(n4510), .A3(n4595), .ZN(n4624) );
  ND3D0 U4237 ( .A1(n4458), .A2(n4051), .A3(n4595), .ZN(n4622) );
  INR3D0 U4238 ( .A1(n4625), .B1(n3273), .B2(n3272), .ZN(n4595) );
  CKND0 U4239 ( .I(n4503), .ZN(n3272) );
  IND2D0 U4240 ( .A1(n4626), .B1(n4627), .ZN(n4503) );
  CKND2D0 U4241 ( .A1(n4501), .A2(n4553), .ZN(n3273) );
  AN3D0 U4242 ( .A1(n4486), .A2(n4433), .A3(n4451), .Z(n4553) );
  CKND2D0 U4243 ( .A1(n4597), .A2(n4593), .ZN(n4451) );
  CKND0 U4244 ( .I(n4628), .ZN(n4597) );
  ND3D0 U4245 ( .A1(n4598), .A2(n4628), .A3(n4593), .ZN(n4433) );
  AN3D0 U4246 ( .A1(n4626), .A2(n4629), .A3(n4627), .Z(n4593) );
  ND3D0 U4247 ( .A1(n4411), .A2(n4062), .A3(n4625), .ZN(n4628) );
  AN3D0 U4248 ( .A1(n4428), .A2(n4060), .A3(n4625), .Z(n4598) );
  IND3D0 U4249 ( .A1(n4629), .B1(n4627), .B2(n4626), .ZN(n4486) );
  ND3D0 U4250 ( .A1(n4557), .A2(n4066), .A3(n4625), .ZN(n4626) );
  AN3D0 U4251 ( .A1(n4630), .A2(n4631), .A3(n4632), .Z(n4627) );
  ND3D0 U4252 ( .A1(n4480), .A2(n4065), .A3(n4625), .ZN(n4629) );
  AN4D0 U4253 ( .A1(n3697), .A2(n4550), .A3(n3696), .A4(n3741), .Z(n4501) );
  IND2D0 U4254 ( .A1(n4633), .B1(n4550), .ZN(n3741) );
  IND2D0 U4255 ( .A1(n4630), .B1(n4632), .ZN(n3696) );
  IND3D0 U4256 ( .A1(n4631), .B1(n4632), .B2(n4630), .ZN(n3697) );
  ND3D0 U4257 ( .A1(n4532), .A2(n4069), .A3(n4625), .ZN(n4630) );
  AN2D0 U4258 ( .A1(n4633), .A2(n4550), .Z(n4632) );
  CKND2D0 U4259 ( .A1(n4625), .A2(n4067), .ZN(n4550) );
  ND3D0 U4260 ( .A1(n4371), .A2(n4510), .A3(n4625), .ZN(n4633) );
  ND3D0 U4261 ( .A1(n4458), .A2(n4070), .A3(n4625), .ZN(n4631) );
  INR2D0 U4262 ( .A1(n3350), .B1(n4575), .ZN(n4625) );
  NR3D0 U4263 ( .A1(n3724), .A2(n4441), .A3(n4440), .ZN(n3350) );
  ND4D0 U4264 ( .A1(n3707), .A2(n4590), .A3(n4474), .A4(n3756), .ZN(n4440) );
  CKND2D0 U4265 ( .A1(n4634), .A2(n4590), .ZN(n3756) );
  CKND2D0 U4266 ( .A1(n4635), .A2(n4636), .ZN(n4474) );
  ND3D0 U4267 ( .A1(n4637), .A2(n4638), .A3(n4639), .ZN(n3707) );
  CKND0 U4268 ( .I(n3706), .ZN(n4441) );
  CKND2D0 U4269 ( .A1(n4640), .A2(n4637), .ZN(n3706) );
  CKND0 U4270 ( .I(n4591), .ZN(n3724) );
  NR2D0 U4271 ( .A1(n3704), .A2(n4442), .ZN(n4591) );
  CKND0 U4272 ( .I(n3755), .ZN(n4442) );
  ND3D0 U4273 ( .A1(n4635), .A2(n4641), .A3(n4642), .ZN(n3755) );
  CKND2D0 U4274 ( .A1(n4446), .A2(n4438), .ZN(n3704) );
  ND3D0 U4275 ( .A1(n4576), .A2(n4643), .A3(n4644), .ZN(n4438) );
  AOI211D0 U4276 ( .A1(n4411), .A2(n4076), .B(n4436), .C(n4077), .ZN(n4644) );
  ND4D0 U4277 ( .A1(n4576), .A2(n4643), .A3(n4411), .A4(n4076), .ZN(n4446) );
  INR3D0 U4278 ( .A1(n4635), .B1(n4642), .B2(n4636), .ZN(n4576) );
  CKND0 U4279 ( .I(n4641), .ZN(n4636) );
  ND3D0 U4280 ( .A1(n4557), .A2(n4083), .A3(n4643), .ZN(n4641) );
  NR3D0 U4281 ( .A1(n4645), .A2(n4074), .A3(n4575), .ZN(n4642) );
  INR3D0 U4282 ( .A1(n4637), .B1(n4639), .B2(n4640), .ZN(n4635) );
  CKND0 U4283 ( .I(n4638), .ZN(n4640) );
  ND3D0 U4284 ( .A1(n4532), .A2(n4082), .A3(n4643), .ZN(n4638) );
  NR3D0 U4285 ( .A1(n4463), .A2(n4004), .A3(n4575), .ZN(n4639) );
  INR2D0 U4286 ( .A1(n4590), .B1(n4634), .ZN(n4637) );
  NR3D0 U4287 ( .A1(n4080), .A2(n4515), .A3(n4575), .ZN(n4634) );
  CKND2D0 U4288 ( .A1(n4643), .A2(n4079), .ZN(n4590) );
  CKND0 U4289 ( .I(n4575), .ZN(n4643) );
  ND3D0 U4290 ( .A1(n4646), .A2(n3314), .A3(n3313), .ZN(n4575) );
  CKND0 U4291 ( .I(n4492), .ZN(n3313) );
  CKND2D0 U4292 ( .A1(n4445), .A2(n4437), .ZN(n4492) );
  ND3D0 U4293 ( .A1(n4581), .A2(n4646), .A3(n4647), .ZN(n4437) );
  AOI211D0 U4294 ( .A1(n4411), .A2(n4097), .B(n4436), .C(n4092), .ZN(n4647) );
  ND4D0 U4295 ( .A1(n4581), .A2(n4646), .A3(n4411), .A4(n4097), .ZN(n4445) );
  AN3D0 U4296 ( .A1(n4648), .A2(n4649), .A3(n4650), .Z(n4581) );
  INR2D0 U4297 ( .A1(n3746), .B1(n4493), .ZN(n3314) );
  ND3D0 U4298 ( .A1(n4548), .A2(n3747), .A3(n4584), .ZN(n4493) );
  AN3D0 U4299 ( .A1(n3709), .A2(n4547), .A3(n3710), .Z(n4584) );
  IND2D0 U4300 ( .A1(n4651), .B1(n4652), .ZN(n3710) );
  IND3D0 U4301 ( .A1(n4653), .B1(n4652), .B2(n4651), .ZN(n3709) );
  CKND2D0 U4302 ( .A1(n4654), .A2(n4547), .ZN(n3747) );
  IND2D0 U4303 ( .A1(n4649), .B1(n4650), .ZN(n4548) );
  IND3D0 U4304 ( .A1(n4648), .B1(n4650), .B2(n4649), .ZN(n3746) );
  ND3D0 U4305 ( .A1(n4557), .A2(n4096), .A3(n4646), .ZN(n4649) );
  AN3D0 U4306 ( .A1(n4651), .A2(n4653), .A3(n4652), .Z(n4650) );
  INR2D0 U4307 ( .A1(n4547), .B1(n4654), .ZN(n4652) );
  NR3D0 U4308 ( .A1(n4099), .A2(n4515), .A3(n4580), .ZN(n4654) );
  CKND2D0 U4309 ( .A1(n4646), .A2(n4098), .ZN(n4547) );
  ND3D0 U4310 ( .A1(n4458), .A2(n4101), .A3(n4646), .ZN(n4653) );
  ND3D0 U4311 ( .A1(n4532), .A2(n4100), .A3(n4646), .ZN(n4651) );
  ND3D0 U4312 ( .A1(n4480), .A2(n4087), .A3(n4646), .ZN(n4648) );
  CKND0 U4313 ( .I(n4580), .ZN(n4646) );
  IND4D0 U4314 ( .A1(n3347), .B1(n3349), .B2(n4655), .B3(n3348), .ZN(n4580) );
  ND3D0 U4315 ( .A1(n4656), .A2(n4655), .A3(n4657), .ZN(n3348) );
  AOI211D0 U4316 ( .A1(n4557), .A2(n4115), .B(n4645), .C(n4114), .ZN(n4657) );
  AN2D0 U4317 ( .A1(n4444), .A2(n4448), .Z(n3349) );
  ND3D0 U4318 ( .A1(n4658), .A2(n4655), .A3(n4659), .ZN(n4448) );
  AOI211D0 U4319 ( .A1(n4411), .A2(n4106), .B(n4436), .C(n4107), .ZN(n4659) );
  ND4D0 U4320 ( .A1(n4658), .A2(n4655), .A3(n4411), .A4(n4106), .ZN(n4444) );
  OA221D0 U4321 ( .A1(n4397), .A2(n4570), .B1(n4114), .B2(n4645), .C(n4656), 
        .Z(n4658) );
  ND4D0 U4322 ( .A1(n4589), .A2(n4543), .A3(n4546), .A4(n4660), .ZN(n3347) );
  AN2D0 U4323 ( .A1(n4586), .A2(n4587), .Z(n4660) );
  IND2D0 U4324 ( .A1(n4661), .B1(n4662), .ZN(n4587) );
  IND3D0 U4325 ( .A1(n4663), .B1(n4662), .B2(n4661), .ZN(n4586) );
  ND4D0 U4326 ( .A1(n4656), .A2(n4655), .A3(n4557), .A4(n4115), .ZN(n4546) );
  AN3D0 U4327 ( .A1(n4661), .A2(n4663), .A3(n4662), .Z(n4656) );
  AN2D0 U4328 ( .A1(n4664), .A2(n4543), .Z(n4662) );
  ND3D0 U4329 ( .A1(n4458), .A2(n4104), .A3(n4655), .ZN(n4663) );
  ND3D0 U4330 ( .A1(n4532), .A2(n4113), .A3(n4655), .ZN(n4661) );
  IND2D0 U4331 ( .A1(n4664), .B1(n4543), .ZN(n4589) );
  CKND2D0 U4332 ( .A1(n4655), .A2(n4112), .ZN(n4543) );
  ND3D0 U4333 ( .A1(n4111), .A2(n4510), .A3(n4655), .ZN(n4664) );
  AN3D0 U4334 ( .A1(n4495), .A2(n4583), .A3(n4494), .Z(n4655) );
  CKND0 U4335 ( .I(n4423), .ZN(n4494) );
  ND4D0 U4336 ( .A1(n4585), .A2(n4150), .A3(n4545), .A4(n4665), .ZN(n4423) );
  OA21D0 U4337 ( .A1(n3937), .A2(n4515), .B(n4588), .Z(n4665) );
  CKND2D0 U4338 ( .A1(n4666), .A2(n4667), .ZN(n4588) );
  IND4D0 U4339 ( .A1(n4668), .B1(n4669), .B2(n4667), .B3(n4670), .ZN(n4545) );
  ND3D0 U4340 ( .A1(n4667), .A2(n4670), .A3(n4668), .ZN(n4585) );
  ND3D0 U4341 ( .A1(n4480), .A2(n4144), .A3(n4671), .ZN(n4583) );
  CKND0 U4342 ( .I(n4645), .ZN(n4480) );
  AN2D0 U4343 ( .A1(n4447), .A2(n4443), .Z(n4495) );
  ND3D0 U4344 ( .A1(n4672), .A2(n4121), .A3(n4411), .ZN(n4443) );
  ND4D0 U4345 ( .A1(n4428), .A2(n4672), .A3(n4119), .A4(n4673), .ZN(n4447) );
  CKND2D0 U4346 ( .A1(n4411), .A2(n4121), .ZN(n4673) );
  CKND0 U4347 ( .I(n4417), .ZN(n4411) );
  OAI221D0 U4348 ( .A1(n4674), .A2(n4675), .B1(n4676), .B2(n3646), .C(n4677), 
        .ZN(n4417) );
  CKND0 U4349 ( .I(n4678), .ZN(n4677) );
  AOI221D0 U4350 ( .A1(n4679), .A2(n4680), .B1(n4681), .B2(n4682), .C(n4683), 
        .ZN(n4676) );
  OAI21D0 U4351 ( .A1(n4684), .A2(n4674), .B(n4685), .ZN(n4682) );
  NR4D0 U4352 ( .A1(n4686), .A2(n4687), .A3(n3680), .A4(n3677), .ZN(n4684) );
  IND2D0 U4353 ( .A1(n3671), .B1(n4688), .ZN(n4679) );
  NR2D0 U4354 ( .A1(n4689), .A2(n4690), .ZN(n4675) );
  OA21D0 U4355 ( .A1(n4146), .A2(n4645), .B(n4671), .Z(n4672) );
  INR4D0 U4356 ( .A1(n4667), .B1(n4668), .B2(n4669), .B3(n4666), .ZN(n4671) );
  CKND0 U4357 ( .I(n4670), .ZN(n4666) );
  CKND2D0 U4358 ( .A1(n4532), .A2(n4151), .ZN(n4670) );
  CKND0 U4359 ( .I(n4537), .ZN(n4532) );
  OAI221D0 U4360 ( .A1(n4691), .A2(n4692), .B1(n4693), .B2(n3648), .C(n4694), 
        .ZN(n4537) );
  AOI221D0 U4361 ( .A1(n4695), .A2(n4696), .B1(n3625), .B2(n4697), .C(n4698), 
        .ZN(n4693) );
  OAI211D0 U4362 ( .A1(n4691), .A2(n4699), .B(n3636), .C(n4700), .ZN(n4697) );
  AOI21D0 U4363 ( .A1(n4681), .A2(n4701), .B(n4702), .ZN(n4700) );
  CKND2D0 U4364 ( .A1(n4703), .A2(n4704), .ZN(n4701) );
  AO21D0 U4365 ( .A1(n4705), .A2(n4706), .B(n4691), .Z(n4704) );
  NR4D0 U4366 ( .A1(n3676), .A2(n3650), .A3(n4707), .A4(n4708), .ZN(n4699) );
  CKND0 U4367 ( .I(n3635), .ZN(n3676) );
  CKND2D0 U4368 ( .A1(n4709), .A2(n4710), .ZN(n4695) );
  INR2D0 U4369 ( .A1(n4711), .B1(n4712), .ZN(n4692) );
  NR2D0 U4370 ( .A1(n4570), .A2(n4456), .ZN(n4669) );
  NR2D0 U4371 ( .A1(n4463), .A2(n4457), .ZN(n4668) );
  CKND2D0 U4372 ( .A1(n4479), .A2(n4510), .ZN(n4667) );
  OAI211D0 U4373 ( .A1(n4713), .A2(n4714), .B(n4715), .C(n4716), .ZN(n4645) );
  AOI21D0 U4374 ( .A1(n4717), .A2(n4718), .B(n4719), .ZN(n4716) );
  OAI21D0 U4375 ( .A1(n4720), .A2(n3639), .B(n3672), .ZN(n4718) );
  NR4D0 U4376 ( .A1(n4721), .A2(n4722), .A3(n3630), .A4(n4707), .ZN(n4714) );
  OAI21D0 U4377 ( .A1(n4723), .A2(n3644), .B(n3632), .ZN(n4722) );
  CKND0 U4378 ( .I(n4717), .ZN(n3644) );
  NR2D0 U4379 ( .A1(n3646), .A2(n3637), .ZN(n4717) );
  NR4D0 U4380 ( .A1(n4724), .A2(n4725), .A3(n4687), .A4(n4726), .ZN(n4723) );
  ND3D0 U4381 ( .A1(n4727), .A2(n4728), .A3(n3611), .ZN(n4724) );
  IIND4D0 U4382 ( .A1(n3619), .A2(n3627), .B1(n4729), .B2(n4730), .ZN(n4721)
         );
  ND3D0 U4383 ( .A1(n4731), .A2(n4732), .A3(n4733), .ZN(n3627) );
  CKND2D0 U4384 ( .A1(n4734), .A2(n4735), .ZN(n3619) );
  CKND0 U4385 ( .I(n4436), .ZN(n4428) );
  OAI221D0 U4386 ( .A1(n4736), .A2(n4737), .B1(n4738), .B2(n3646), .C(n4739), 
        .ZN(n4436) );
  CKND0 U4387 ( .I(n4689), .ZN(n4739) );
  OAI21D0 U4388 ( .A1(n3663), .A2(n3648), .B(n4734), .ZN(n4689) );
  CKND0 U4389 ( .I(n3662), .ZN(n4734) );
  CKND2D0 U4390 ( .A1(n4740), .A2(n4741), .ZN(n3662) );
  AN2D0 U4391 ( .A1(n4732), .A2(n4742), .Z(n3663) );
  CKND2D0 U4392 ( .A1(n3617), .A2(n3625), .ZN(n3646) );
  CKND0 U4393 ( .I(n3648), .ZN(n3617) );
  AOI221D0 U4394 ( .A1(n4681), .A2(n3677), .B1(n4743), .B2(n4744), .C(n3671), 
        .ZN(n4738) );
  CKND2D0 U4395 ( .A1(n4745), .A2(n4746), .ZN(n3671) );
  IND4D0 U4396 ( .A1(n4683), .B1(n4685), .B2(n4688), .B3(n4747), .ZN(n4743) );
  NR3D0 U4397 ( .A1(n3680), .A2(n4686), .A3(n4687), .ZN(n4747) );
  INR4D0 U4398 ( .A1(n3326), .B1(n4707), .B2(n4702), .B3(n4719), .ZN(n4688) );
  AN2D0 U4399 ( .A1(n4748), .A2(n4749), .Z(n4685) );
  CKND2D0 U4400 ( .A1(n4750), .A2(n4751), .ZN(n4683) );
  CKND2D0 U4401 ( .A1(n4752), .A2(n4753), .ZN(n3677) );
  NR2D0 U4402 ( .A1(n4690), .A2(n4678), .ZN(n4737) );
  CKND2D0 U4403 ( .A1(n4735), .A2(n4754), .ZN(n4678) );
  AO21D0 U4404 ( .A1(n4731), .A2(n4755), .B(n3648), .Z(n4754) );
  OA21D0 U4405 ( .A1(n4756), .A2(n4757), .B(n4758), .Z(n4735) );
  OAI211D0 U4406 ( .A1(n4729), .A2(n3648), .B(n4730), .C(n4715), .ZN(n4690) );
  OA211D0 U4407 ( .A1(n3665), .A2(n3648), .B(n3655), .C(n3658), .Z(n4715) );
  AN2D0 U4408 ( .A1(n4759), .A2(n4760), .Z(n3665) );
  AN2D0 U4409 ( .A1(n3296), .A2(n4761), .Z(n4730) );
  AN4D0 U4410 ( .A1(n3660), .A2(n4762), .A3(n3613), .A4(n4763), .Z(n3296) );
  NR2D0 U4411 ( .A1(n4764), .A2(n3620), .ZN(n4763) );
  AN4D0 U4412 ( .A1(n4765), .A2(n4766), .A3(n4767), .A4(n4768), .Z(n4729) );
  CKND0 U4413 ( .I(n4515), .ZN(n4510) );
  OAI221D0 U4414 ( .A1(n4769), .A2(n4770), .B1(n4771), .B2(n3648), .C(n4772), 
        .ZN(n4515) );
  AOI221D0 U4415 ( .A1(n4773), .A2(n4774), .B1(n3625), .B2(n4775), .C(n4776), 
        .ZN(n4771) );
  OAI221D0 U4416 ( .A1(n4769), .A2(n4777), .B1(n4778), .B2(n3637), .C(n3682), 
        .ZN(n4775) );
  AOI221D0 U4417 ( .A1(n3651), .A2(n3679), .B1(n4779), .B2(n4774), .C(n4780), 
        .ZN(n4778) );
  ND4D0 U4418 ( .A1(n4781), .A2(n4703), .A3(n4782), .A4(n4706), .ZN(n4779) );
  NR2D0 U4419 ( .A1(n4783), .A2(n3652), .ZN(n4782) );
  NR2D0 U4420 ( .A1(n3649), .A2(n4784), .ZN(n4777) );
  CKND0 U4421 ( .I(n4785), .ZN(n3649) );
  CKND2D0 U4422 ( .A1(n4786), .A2(n4710), .ZN(n4773) );
  INR2D0 U4423 ( .A1(n4787), .B1(n4788), .ZN(n4710) );
  NR3D0 U4424 ( .A1(n4789), .A2(n4790), .A3(n4712), .ZN(n4770) );
  ND3D0 U4425 ( .A1(n3654), .A2(n4762), .A3(n4791), .ZN(n4712) );
  CKND0 U4426 ( .I(n4463), .ZN(n4458) );
  OAI221D0 U4427 ( .A1(n4792), .A2(n4793), .B1(n4794), .B2(n3648), .C(n4795), 
        .ZN(n4463) );
  AOI221D0 U4428 ( .A1(n4796), .A2(n4797), .B1(n3625), .B2(n4798), .C(n4788), 
        .ZN(n4794) );
  CKND2D0 U4429 ( .A1(n3629), .A2(n3623), .ZN(n4788) );
  ND4D0 U4430 ( .A1(n4799), .A2(n3635), .A3(n4800), .A4(n3633), .ZN(n4798) );
  OAI21D0 U4431 ( .A1(n4801), .A2(n3678), .B(n4681), .ZN(n4800) );
  NR2D0 U4432 ( .A1(n3637), .A2(n3639), .ZN(n4681) );
  AOI21D0 U4433 ( .A1(n4703), .A2(n4705), .B(n4792), .ZN(n4801) );
  INR3D0 U4434 ( .A1(n4802), .B1(n3679), .B2(n3652), .ZN(n4705) );
  ND4D0 U4435 ( .A1(n4720), .A2(n3611), .A3(n4803), .A4(n4728), .ZN(n3652) );
  AN2D0 U4436 ( .A1(n4804), .A2(n4805), .Z(n4803) );
  CKND0 U4437 ( .I(n3680), .ZN(n4720) );
  OAI31D0 U4438 ( .A1(n4806), .A2(n4708), .A3(n4807), .B(n4797), .ZN(n4799) );
  IND3D0 U4439 ( .A1(n3653), .B1(n4808), .B2(n3673), .ZN(n4708) );
  ND3D0 U4440 ( .A1(n3672), .A2(n4809), .A3(n3325), .ZN(n3653) );
  ND3D0 U4441 ( .A1(n4785), .A2(n3682), .A3(n3636), .ZN(n4806) );
  ND3D0 U4442 ( .A1(n4709), .A2(n4787), .A3(n4786), .ZN(n4796) );
  CKND0 U4443 ( .I(n4698), .ZN(n4786) );
  CKND2D0 U4444 ( .A1(n3621), .A2(n3622), .ZN(n4698) );
  AN3D0 U4445 ( .A1(n4810), .A2(n4811), .A3(n3647), .Z(n4787) );
  AN3D0 U4446 ( .A1(n4812), .A2(n4813), .A3(n4814), .Z(n3647) );
  CKND0 U4447 ( .I(n4815), .ZN(n4812) );
  CKND0 U4448 ( .I(n4776), .ZN(n4709) );
  CKND2D0 U4449 ( .A1(n3668), .A2(n3667), .ZN(n4776) );
  NR2D0 U4450 ( .A1(n4816), .A2(n4817), .ZN(n4793) );
  CKND0 U4451 ( .I(n4570), .ZN(n4557) );
  OAI221D0 U4452 ( .A1(n4818), .A2(n4819), .B1(n4820), .B2(n3648), .C(n3642), 
        .ZN(n4570) );
  CKND0 U4453 ( .I(n4817), .ZN(n3642) );
  CKND2D0 U4454 ( .A1(n4762), .A2(n4821), .ZN(n4817) );
  ND4D0 U4455 ( .A1(n4822), .A2(n4823), .A3(n4824), .A4(n4825), .ZN(n4762) );
  ND3D0 U4456 ( .A1(n4826), .A2(n4827), .A3(n4828), .ZN(n3648) );
  AOI221D0 U4457 ( .A1(n4829), .A2(n4830), .B1(n3625), .B2(n4831), .C(n4815), 
        .ZN(n4820) );
  CKND2D0 U4458 ( .A1(n4767), .A2(n4768), .ZN(n4815) );
  OAI221D0 U4459 ( .A1(n4818), .A2(n4832), .B1(n4833), .B2(n3637), .C(n4785), 
        .ZN(n4831) );
  OAI21D0 U4460 ( .A1(n4834), .A2(n4835), .B(n4836), .ZN(n3637) );
  AOI22D0 U4461 ( .A1(n4736), .A2(n4326), .B1(n4674), .B2(n4076), .ZN(n4834)
         );
  AOI221D0 U4462 ( .A1(n4837), .A2(n4830), .B1(n3651), .B2(n4838), .C(n4783), 
        .ZN(n4833) );
  CKND0 U4463 ( .I(n4809), .ZN(n4783) );
  CKND2D0 U4464 ( .A1(n4804), .A2(n4805), .ZN(n4838) );
  CKND0 U4465 ( .I(n3639), .ZN(n3651) );
  OAI21D0 U4466 ( .A1(n4839), .A2(n4840), .B(n4841), .ZN(n3639) );
  AOI22D0 U4467 ( .A1(n4736), .A2(n4310), .B1(n4674), .B2(n4097), .ZN(n4839)
         );
  IND4D0 U4468 ( .A1(n3679), .B1(n3638), .B2(n4781), .B3(n4842), .ZN(n4837) );
  NR2D0 U4469 ( .A1(n4780), .A2(n3680), .ZN(n4842) );
  CKND2D0 U4470 ( .A1(n4843), .A2(n3610), .ZN(n3680) );
  CKND0 U4471 ( .I(n3673), .ZN(n4780) );
  AN4D0 U4472 ( .A1(n3325), .A2(n4844), .A3(n3672), .A4(n4802), .Z(n4781) );
  AN4D0 U4473 ( .A1(n4703), .A2(n4706), .A3(n3611), .A4(n4728), .Z(n3638) );
  CKND0 U4474 ( .I(n3678), .ZN(n4706) );
  CKND2D0 U4475 ( .A1(n4845), .A2(n4846), .ZN(n3678) );
  AN2D0 U4476 ( .A1(n4847), .A2(n4848), .Z(n4703) );
  OAI21D0 U4477 ( .A1(n4774), .A2(n3937), .B(n4849), .ZN(n3679) );
  INR2D0 U4478 ( .A1(n3682), .B1(n4784), .ZN(n4832) );
  IND2D0 U4479 ( .A1(n4807), .B1(n3633), .ZN(n4784) );
  ND3D0 U4480 ( .A1(n3632), .A2(n4850), .A3(n4851), .ZN(n4807) );
  AN3D0 U4481 ( .A1(n4852), .A2(n4853), .A3(n4854), .Z(n3625) );
  AOI211D0 U4482 ( .A1(n4855), .A2(n4856), .B(n4857), .C(n4858), .ZN(n4854) );
  OAI22D0 U4483 ( .A1(n4302), .A2(n4680), .B1(n4043), .B2(n4744), .ZN(n4856)
         );
  IND3D0 U4484 ( .A1(n3300), .B1(n4765), .B2(n4813), .ZN(n4829) );
  INR2D0 U4485 ( .A1(n4795), .B1(n4816), .ZN(n4819) );
  CKND2D0 U4486 ( .A1(n4694), .A2(n4711), .ZN(n4816) );
  INR2D0 U4487 ( .A1(n4772), .B1(n4790), .ZN(n4711) );
  ND3D0 U4488 ( .A1(n4859), .A2(n4860), .A3(n3641), .ZN(n4790) );
  AN2D0 U4489 ( .A1(n3294), .A2(n4861), .Z(n3641) );
  AN3D0 U4490 ( .A1(n3655), .A2(n4758), .A3(n4741), .Z(n3294) );
  ND3D0 U4491 ( .A1(n4828), .A2(n4824), .A3(n4862), .ZN(n4741) );
  AOI211D0 U4492 ( .A1(n4674), .A2(n3946), .B(n4744), .C(n3373), .ZN(n4862) );
  ND4D0 U4493 ( .A1(n4828), .A2(n4824), .A3(n4674), .A4(n3946), .ZN(n4758) );
  OA211D0 U4494 ( .A1(n4863), .A2(n4864), .B(n4825), .C(n4823), .Z(n4828) );
  CKND0 U4495 ( .I(n4865), .ZN(n4825) );
  AOI21D0 U4496 ( .A1(n4713), .A2(n4014), .B(n4822), .ZN(n4863) );
  ND4D0 U4497 ( .A1(n4824), .A2(n4713), .A3(n4823), .A4(n4866), .ZN(n3655) );
  NR3D0 U4498 ( .A1(n3372), .A2(n4822), .A3(n4865), .ZN(n4866) );
  INR2D0 U4499 ( .A1(n4016), .B1(n4830), .ZN(n4822) );
  AN2D0 U4500 ( .A1(n3660), .A2(n3659), .Z(n4772) );
  OR2D0 U4501 ( .A1(n4867), .A2(n4764), .Z(n3660) );
  CKND0 U4502 ( .I(n4859), .ZN(n4764) );
  CKND0 U4503 ( .I(n4789), .ZN(n4694) );
  CKND2D0 U4504 ( .A1(n3613), .A2(n3614), .ZN(n4789) );
  IND3D0 U4505 ( .A1(n4868), .B1(n4867), .B2(n4859), .ZN(n3613) );
  INR2D0 U4506 ( .A1(n3615), .B1(n3620), .ZN(n4795) );
  CKND0 U4507 ( .I(n3654), .ZN(n3620) );
  CKND2D0 U4508 ( .A1(n4865), .A2(n4823), .ZN(n3654) );
  AN3D0 U4509 ( .A1(n4868), .A2(n4859), .A3(n4867), .Z(n4823) );
  IND3D0 U4510 ( .A1(n3894), .B1(n4769), .B2(n4824), .ZN(n4867) );
  CKND2D0 U4511 ( .A1(n4824), .A2(n3893), .ZN(n4859) );
  ND3D0 U4512 ( .A1(n4691), .A2(n4019), .A3(n4824), .ZN(n4868) );
  CKND0 U4513 ( .I(n4864), .ZN(n4824) );
  NR3D0 U4514 ( .A1(n4797), .A2(n4011), .A3(n4864), .ZN(n4865) );
  CKND2D0 U4515 ( .A1(n3295), .A2(n4869), .ZN(n4864) );
  AN2D0 U4516 ( .A1(n4761), .A2(n4861), .Z(n3295) );
  OA211D0 U4517 ( .A1(n4756), .A2(n4757), .B(n3658), .C(n4740), .Z(n4861) );
  IND3D0 U4518 ( .A1(n4827), .B1(n4757), .B2(n4826), .ZN(n4740) );
  CKND0 U4519 ( .I(n4756), .ZN(n4826) );
  ND3D0 U4520 ( .A1(n4736), .A2(n4028), .A3(n4869), .ZN(n4827) );
  IND3D0 U4521 ( .A1(n4870), .B1(n4871), .B2(n4872), .ZN(n3658) );
  ND3D0 U4522 ( .A1(n4674), .A2(n4034), .A3(n4869), .ZN(n4757) );
  ND3D0 U4523 ( .A1(n4870), .A2(n4872), .A3(n4871), .ZN(n4756) );
  ND3D0 U4524 ( .A1(n4713), .A2(n4029), .A3(n4869), .ZN(n4870) );
  AN4D0 U4525 ( .A1(n4791), .A2(n4860), .A3(n3614), .A4(n3659), .Z(n4761) );
  IND2D0 U4526 ( .A1(n4873), .B1(n4860), .ZN(n3659) );
  IND2D0 U4527 ( .A1(n4874), .B1(n4875), .ZN(n3614) );
  AN2D0 U4528 ( .A1(n4821), .A2(n3615), .Z(n4791) );
  IND2D0 U4529 ( .A1(n4872), .B1(n4871), .ZN(n4821) );
  AN3D0 U4530 ( .A1(n4874), .A2(n4876), .A3(n4875), .Z(n4871) );
  ND3D0 U4531 ( .A1(n4818), .A2(n4033), .A3(n4869), .ZN(n4872) );
  IND3D0 U4532 ( .A1(n4876), .B1(n4875), .B2(n4874), .ZN(n3615) );
  ND3D0 U4533 ( .A1(n4691), .A2(n4037), .A3(n4869), .ZN(n4874) );
  AN2D0 U4534 ( .A1(n4873), .A2(n4860), .Z(n4875) );
  CKND2D0 U4535 ( .A1(n4869), .A2(n4035), .ZN(n4860) );
  ND3D0 U4536 ( .A1(n4352), .A2(n4769), .A3(n4869), .ZN(n4873) );
  ND3D0 U4537 ( .A1(n4792), .A2(n4038), .A3(n4869), .ZN(n4876) );
  INR2D0 U4538 ( .A1(n4855), .B1(n3298), .ZN(n4869) );
  ND3D0 U4539 ( .A1(n4765), .A2(n4767), .A3(n4813), .ZN(n3298) );
  AN2D0 U4540 ( .A1(n4733), .A2(n4760), .Z(n4813) );
  IND3D0 U4541 ( .A1(n4877), .B1(n4878), .B2(n4879), .ZN(n4760) );
  AN2D0 U4542 ( .A1(n4755), .A2(n4742), .Z(n4733) );
  ND3D0 U4543 ( .A1(n4852), .A2(n4855), .A3(n4880), .ZN(n4742) );
  AOI211D0 U4544 ( .A1(n4674), .A2(n4042), .B(n4744), .C(n4043), .ZN(n4880) );
  ND4D0 U4545 ( .A1(n4852), .A2(n4855), .A3(n4674), .A4(n4042), .ZN(n4755) );
  AN3D0 U4546 ( .A1(n4877), .A2(n4879), .A3(n4878), .Z(n4852) );
  ND3D0 U4547 ( .A1(n4713), .A2(n4047), .A3(n4855), .ZN(n4877) );
  IND2D0 U4548 ( .A1(n4879), .B1(n4878), .ZN(n4767) );
  AN3D0 U4549 ( .A1(n4881), .A2(n4882), .A3(n4883), .Z(n4878) );
  ND3D0 U4550 ( .A1(n4818), .A2(n4053), .A3(n4855), .ZN(n4879) );
  AN4D0 U4551 ( .A1(n3629), .A2(n4810), .A3(n3621), .A4(n3668), .Z(n4765) );
  IND2D0 U4552 ( .A1(n4884), .B1(n4810), .ZN(n3668) );
  IND2D0 U4553 ( .A1(n4881), .B1(n4883), .ZN(n3621) );
  IND3D0 U4554 ( .A1(n4882), .B1(n4883), .B2(n4881), .ZN(n3629) );
  ND3D0 U4555 ( .A1(n4691), .A2(n4052), .A3(n4855), .ZN(n4881) );
  AN2D0 U4556 ( .A1(n4884), .A2(n4810), .Z(n4883) );
  CKND2D0 U4557 ( .A1(n4855), .A2(n4049), .ZN(n4810) );
  ND3D0 U4558 ( .A1(n4361), .A2(n4769), .A3(n4855), .ZN(n4884) );
  ND3D0 U4559 ( .A1(n4792), .A2(n4051), .A3(n4855), .ZN(n4882) );
  INR3D0 U4560 ( .A1(n4885), .B1(n3300), .B2(n3299), .ZN(n4855) );
  CKND0 U4561 ( .I(n4768), .ZN(n3299) );
  IND2D0 U4562 ( .A1(n4886), .B1(n4887), .ZN(n4768) );
  CKND2D0 U4563 ( .A1(n4766), .A2(n4814), .ZN(n3300) );
  AN3D0 U4564 ( .A1(n4759), .A2(n4732), .A3(n4731), .Z(n4814) );
  CKND2D0 U4565 ( .A1(n4857), .A2(n4853), .ZN(n4731) );
  CKND0 U4566 ( .I(n4888), .ZN(n4857) );
  ND3D0 U4567 ( .A1(n4858), .A2(n4888), .A3(n4853), .ZN(n4732) );
  AN3D0 U4568 ( .A1(n4886), .A2(n4889), .A3(n4887), .Z(n4853) );
  ND3D0 U4569 ( .A1(n4674), .A2(n4062), .A3(n4885), .ZN(n4888) );
  AN3D0 U4570 ( .A1(n4736), .A2(n4060), .A3(n4885), .Z(n4858) );
  IND3D0 U4571 ( .A1(n4889), .B1(n4887), .B2(n4886), .ZN(n4759) );
  ND3D0 U4572 ( .A1(n4818), .A2(n4066), .A3(n4885), .ZN(n4886) );
  AN3D0 U4573 ( .A1(n4890), .A2(n4891), .A3(n4892), .Z(n4887) );
  ND3D0 U4574 ( .A1(n4713), .A2(n4065), .A3(n4885), .ZN(n4889) );
  AN4D0 U4575 ( .A1(n3623), .A2(n4811), .A3(n3622), .A4(n3667), .Z(n4766) );
  IND2D0 U4576 ( .A1(n4893), .B1(n4811), .ZN(n3667) );
  IND2D0 U4577 ( .A1(n4890), .B1(n4892), .ZN(n3622) );
  IND3D0 U4578 ( .A1(n4891), .B1(n4892), .B2(n4890), .ZN(n3623) );
  ND3D0 U4579 ( .A1(n4691), .A2(n4069), .A3(n4885), .ZN(n4890) );
  AN2D0 U4580 ( .A1(n4893), .A2(n4811), .Z(n4892) );
  CKND2D0 U4581 ( .A1(n4885), .A2(n4067), .ZN(n4811) );
  ND3D0 U4582 ( .A1(n4371), .A2(n4769), .A3(n4885), .ZN(n4893) );
  ND3D0 U4583 ( .A1(n4792), .A2(n4070), .A3(n4885), .ZN(n4891) );
  INR2D0 U4584 ( .A1(n3612), .B1(n4835), .ZN(n4885) );
  NR3D0 U4585 ( .A1(n3650), .A2(n4702), .A3(n4707), .ZN(n3612) );
  ND4D0 U4586 ( .A1(n3633), .A2(n4850), .A3(n4785), .A4(n3682), .ZN(n4707) );
  CKND2D0 U4587 ( .A1(n4894), .A2(n4850), .ZN(n3682) );
  CKND2D0 U4588 ( .A1(n4895), .A2(n4896), .ZN(n4785) );
  ND3D0 U4589 ( .A1(n4897), .A2(n4898), .A3(n4899), .ZN(n3633) );
  CKND0 U4590 ( .I(n3632), .ZN(n4702) );
  CKND2D0 U4591 ( .A1(n4900), .A2(n4897), .ZN(n3632) );
  CKND0 U4592 ( .I(n4851), .ZN(n3650) );
  NR2D0 U4593 ( .A1(n3630), .A2(n4719), .ZN(n4851) );
  CKND0 U4594 ( .I(n3681), .ZN(n4719) );
  ND3D0 U4595 ( .A1(n4895), .A2(n4901), .A3(n4902), .ZN(n3681) );
  CKND2D0 U4596 ( .A1(n4751), .A2(n4746), .ZN(n3630) );
  ND3D0 U4597 ( .A1(n4836), .A2(n4903), .A3(n4904), .ZN(n4746) );
  AOI211D0 U4598 ( .A1(n4674), .A2(n4076), .B(n4744), .C(n4077), .ZN(n4904) );
  ND4D0 U4599 ( .A1(n4836), .A2(n4903), .A3(n4674), .A4(n4076), .ZN(n4751) );
  INR3D0 U4600 ( .A1(n4895), .B1(n4902), .B2(n4896), .ZN(n4836) );
  CKND0 U4601 ( .I(n4901), .ZN(n4896) );
  ND3D0 U4602 ( .A1(n4818), .A2(n4083), .A3(n4903), .ZN(n4901) );
  NR3D0 U4603 ( .A1(n4905), .A2(n4074), .A3(n4835), .ZN(n4902) );
  INR3D0 U4604 ( .A1(n4897), .B1(n4899), .B2(n4900), .ZN(n4895) );
  CKND0 U4605 ( .I(n4898), .ZN(n4900) );
  ND3D0 U4606 ( .A1(n4691), .A2(n4082), .A3(n4903), .ZN(n4898) );
  NR3D0 U4607 ( .A1(n4797), .A2(n4004), .A3(n4835), .ZN(n4899) );
  INR2D0 U4608 ( .A1(n4850), .B1(n4894), .ZN(n4897) );
  NR3D0 U4609 ( .A1(n4080), .A2(n4774), .A3(n4835), .ZN(n4894) );
  CKND2D0 U4610 ( .A1(n4903), .A2(n4079), .ZN(n4850) );
  CKND0 U4611 ( .I(n4835), .ZN(n4903) );
  ND3D0 U4612 ( .A1(n4906), .A2(n3326), .A3(n3325), .ZN(n4835) );
  CKND0 U4613 ( .I(n4725), .ZN(n3325) );
  CKND2D0 U4614 ( .A1(n4750), .A2(n4745), .ZN(n4725) );
  ND3D0 U4615 ( .A1(n4841), .A2(n4906), .A3(n4907), .ZN(n4745) );
  AOI211D0 U4616 ( .A1(n4674), .A2(n4097), .B(n4744), .C(n4092), .ZN(n4907) );
  ND4D0 U4617 ( .A1(n4841), .A2(n4906), .A3(n4674), .A4(n4097), .ZN(n4750) );
  AN3D0 U4618 ( .A1(n4908), .A2(n4909), .A3(n4910), .Z(n4841) );
  INR2D0 U4619 ( .A1(n3672), .B1(n4726), .ZN(n3326) );
  ND3D0 U4620 ( .A1(n4809), .A2(n3673), .A3(n4844), .ZN(n4726) );
  AN3D0 U4621 ( .A1(n3635), .A2(n4808), .A3(n3636), .Z(n4844) );
  IND2D0 U4622 ( .A1(n4911), .B1(n4912), .ZN(n3636) );
  IND3D0 U4623 ( .A1(n4913), .B1(n4912), .B2(n4911), .ZN(n3635) );
  CKND2D0 U4624 ( .A1(n4914), .A2(n4808), .ZN(n3673) );
  IND2D0 U4625 ( .A1(n4909), .B1(n4910), .ZN(n4809) );
  IND3D0 U4626 ( .A1(n4908), .B1(n4910), .B2(n4909), .ZN(n3672) );
  ND3D0 U4627 ( .A1(n4818), .A2(n4096), .A3(n4906), .ZN(n4909) );
  AN3D0 U4628 ( .A1(n4911), .A2(n4913), .A3(n4912), .Z(n4910) );
  INR2D0 U4629 ( .A1(n4808), .B1(n4914), .ZN(n4912) );
  NR3D0 U4630 ( .A1(n4099), .A2(n4774), .A3(n4840), .ZN(n4914) );
  CKND2D0 U4631 ( .A1(n4906), .A2(n4098), .ZN(n4808) );
  ND3D0 U4632 ( .A1(n4792), .A2(n4101), .A3(n4906), .ZN(n4913) );
  ND3D0 U4633 ( .A1(n4691), .A2(n4100), .A3(n4906), .ZN(n4911) );
  ND3D0 U4634 ( .A1(n4713), .A2(n4087), .A3(n4906), .ZN(n4908) );
  CKND0 U4635 ( .I(n4840), .ZN(n4906) );
  ND4D0 U4636 ( .A1(n3609), .A2(n3611), .A3(n4915), .A4(n3610), .ZN(n4840) );
  ND3D0 U4637 ( .A1(n4916), .A2(n4915), .A3(n4917), .ZN(n3610) );
  AOI211D0 U4638 ( .A1(n4818), .A2(n4115), .B(n4905), .C(n4114), .ZN(n4917) );
  AN2D0 U4639 ( .A1(n4749), .A2(n4753), .Z(n3611) );
  ND3D0 U4640 ( .A1(n4918), .A2(n4915), .A3(n4919), .ZN(n4753) );
  AOI211D0 U4641 ( .A1(n4674), .A2(n4106), .B(n4744), .C(n4107), .ZN(n4919) );
  ND4D0 U4642 ( .A1(n4918), .A2(n4915), .A3(n4674), .A4(n4106), .ZN(n4749) );
  OA221D0 U4643 ( .A1(n4397), .A2(n4830), .B1(n4114), .B2(n4905), .C(n4916), 
        .Z(n4918) );
  CKND0 U4644 ( .I(n4687), .ZN(n3609) );
  ND4D0 U4645 ( .A1(n4849), .A2(n4802), .A3(n4805), .A4(n4920), .ZN(n4687) );
  AN2D0 U4646 ( .A1(n4846), .A2(n4847), .Z(n4920) );
  IND2D0 U4647 ( .A1(n4921), .B1(n4922), .ZN(n4847) );
  IND3D0 U4648 ( .A1(n4923), .B1(n4922), .B2(n4921), .ZN(n4846) );
  ND4D0 U4649 ( .A1(n4916), .A2(n4915), .A3(n4818), .A4(n4115), .ZN(n4805) );
  AN3D0 U4650 ( .A1(n4921), .A2(n4923), .A3(n4922), .Z(n4916) );
  AN2D0 U4651 ( .A1(n4924), .A2(n4802), .Z(n4922) );
  ND3D0 U4652 ( .A1(n4792), .A2(n4104), .A3(n4915), .ZN(n4923) );
  ND3D0 U4653 ( .A1(n4691), .A2(n4113), .A3(n4915), .ZN(n4921) );
  IND2D0 U4654 ( .A1(n4924), .B1(n4802), .ZN(n4849) );
  CKND2D0 U4655 ( .A1(n4915), .A2(n4112), .ZN(n4802) );
  ND3D0 U4656 ( .A1(n4111), .A2(n4769), .A3(n4915), .ZN(n4924) );
  AN3D0 U4657 ( .A1(n4728), .A2(n4843), .A3(n4727), .Z(n4915) );
  CKND0 U4658 ( .I(n4686), .ZN(n4727) );
  ND4D0 U4659 ( .A1(n4845), .A2(n4150), .A3(n4804), .A4(n4925), .ZN(n4686) );
  OA21D0 U4660 ( .A1(n3937), .A2(n4774), .B(n4848), .Z(n4925) );
  CKND2D0 U4661 ( .A1(n4926), .A2(n4927), .ZN(n4848) );
  IND4D0 U4662 ( .A1(n4928), .B1(n4929), .B2(n4927), .B3(n4930), .ZN(n4804) );
  ND3D0 U4663 ( .A1(n4927), .A2(n4930), .A3(n4928), .ZN(n4845) );
  ND3D0 U4664 ( .A1(n4713), .A2(n4144), .A3(n4931), .ZN(n4843) );
  CKND0 U4665 ( .I(n4905), .ZN(n4713) );
  AN2D0 U4666 ( .A1(n4752), .A2(n4748), .Z(n4728) );
  ND3D0 U4667 ( .A1(n4932), .A2(n4121), .A3(n4674), .ZN(n4748) );
  ND4D0 U4668 ( .A1(n4736), .A2(n4932), .A3(n4119), .A4(n4933), .ZN(n4752) );
  CKND2D0 U4669 ( .A1(n4674), .A2(n4121), .ZN(n4933) );
  CKND0 U4670 ( .I(n4680), .ZN(n4674) );
  OAI221D0 U4671 ( .A1(n4934), .A2(n4935), .B1(n4936), .B2(n3525), .C(n4937), 
        .ZN(n4680) );
  CKND0 U4672 ( .I(n4938), .ZN(n4937) );
  AOI221D0 U4673 ( .A1(n4939), .A2(n4940), .B1(n3531), .B2(n4941), .C(n4942), 
        .ZN(n4936) );
  OAI211D0 U4674 ( .A1(n4943), .A2(n3556), .B(n4944), .C(n4945), .ZN(n4939) );
  CKND0 U4675 ( .I(n4946), .ZN(n4944) );
  NR2D0 U4676 ( .A1(n4947), .A2(n4948), .ZN(n4935) );
  OA21D0 U4677 ( .A1(n4146), .A2(n4905), .B(n4931), .Z(n4932) );
  INR4D0 U4678 ( .A1(n4927), .B1(n4928), .B2(n4929), .B3(n4926), .ZN(n4931) );
  CKND0 U4679 ( .I(n4930), .ZN(n4926) );
  CKND2D0 U4680 ( .A1(n4691), .A2(n4151), .ZN(n4930) );
  CKND0 U4681 ( .I(n4696), .ZN(n4691) );
  OAI221D0 U4682 ( .A1(n4949), .A2(n4950), .B1(n4951), .B2(n3527), .C(n4952), 
        .ZN(n4696) );
  CKND0 U4683 ( .I(n4953), .ZN(n4952) );
  AOI221D0 U4684 ( .A1(n4954), .A2(n4955), .B1(n3550), .B2(n4956), .C(n4957), 
        .ZN(n4951) );
  OAI211D0 U4685 ( .A1(n4949), .A2(n4958), .B(n4959), .C(n4960), .ZN(n4956) );
  AOI21D0 U4686 ( .A1(n3531), .A2(n4961), .B(n4962), .ZN(n4960) );
  IND2D0 U4687 ( .A1(n4963), .B1(n4964), .ZN(n4961) );
  OAI21D0 U4688 ( .A1(n4965), .A2(n4966), .B(n4955), .ZN(n4964) );
  NR4D0 U4689 ( .A1(n3587), .A2(n3534), .A3(n4967), .A4(n4968), .ZN(n4958) );
  CKND2D0 U4690 ( .A1(n4969), .A2(n4970), .ZN(n4954) );
  NR2D0 U4691 ( .A1(n4971), .A2(n4972), .ZN(n4950) );
  NR2D0 U4692 ( .A1(n4830), .A2(n4456), .ZN(n4929) );
  NR2D0 U4693 ( .A1(n4797), .A2(n4457), .ZN(n4928) );
  CKND2D0 U4694 ( .A1(n4479), .A2(n4769), .ZN(n4927) );
  OAI221D0 U4695 ( .A1(n4973), .A2(n3525), .B1(n4974), .B2(n4975), .C(n4976), 
        .ZN(n4905) );
  NR4D0 U4696 ( .A1(n4977), .A2(n3544), .A3(n3552), .A4(n4978), .ZN(n4975) );
  ND3D0 U4697 ( .A1(n4979), .A2(n4980), .A3(n4981), .ZN(n3552) );
  CKND2D0 U4698 ( .A1(n3565), .A2(n4982), .ZN(n3544) );
  IND4D0 U4699 ( .A1(n4967), .B1(n4983), .B2(n3557), .B3(n4959), .ZN(n4977) );
  AOI221D0 U4700 ( .A1(n4984), .A2(n4985), .B1(n3531), .B2(n3594), .C(n4986), 
        .ZN(n4973) );
  ND4D0 U4701 ( .A1(n4987), .A2(n3311), .A3(n4988), .A4(n4989), .ZN(n4984) );
  NR2D0 U4702 ( .A1(n3563), .A2(n4990), .ZN(n4989) );
  CKND0 U4703 ( .I(n4744), .ZN(n4736) );
  OAI221D0 U4704 ( .A1(n4991), .A2(n4992), .B1(n4993), .B2(n3525), .C(n4994), 
        .ZN(n4744) );
  CKND0 U4705 ( .I(n4947), .ZN(n4994) );
  OAI21D0 U4706 ( .A1(n3577), .A2(n3527), .B(n3565), .ZN(n4947) );
  AN2D0 U4707 ( .A1(n4995), .A2(n4996), .Z(n3565) );
  AN2D0 U4708 ( .A1(n4980), .A2(n4997), .Z(n3577) );
  CKND2D0 U4709 ( .A1(n3542), .A2(n3550), .ZN(n3525) );
  CKND0 U4710 ( .I(n3527), .ZN(n3542) );
  AOI21D0 U4711 ( .A1(n4998), .A2(n4999), .B(n4946), .ZN(n4993) );
  OAI211D0 U4712 ( .A1(n5000), .A2(n3556), .B(n3584), .C(n3580), .ZN(n4946) );
  NR2D0 U4713 ( .A1(n3596), .A2(n3595), .ZN(n5000) );
  CKND0 U4714 ( .I(n5001), .ZN(n3595) );
  CKND0 U4715 ( .I(n5002), .ZN(n3596) );
  IIND4D0 U4716 ( .A1(n4941), .A2(n4942), .B1(n4943), .B2(n4945), .ZN(n4998)
         );
  INR4D0 U4717 ( .A1(n3311), .B1(n4986), .B2(n4967), .B3(n3562), .ZN(n4945) );
  CKND2D0 U4718 ( .A1(n3582), .A2(n5003), .ZN(n4986) );
  NR2D0 U4719 ( .A1(n4990), .A2(n3594), .ZN(n4943) );
  IND4D0 U4720 ( .A1(n5004), .B1(n3338), .B2(n5005), .B3(n5006), .ZN(n4990) );
  CKND2D0 U4721 ( .A1(n5007), .A2(n5008), .ZN(n4942) );
  CKND2D0 U4722 ( .A1(n5009), .A2(n5010), .ZN(n4941) );
  NR2D0 U4723 ( .A1(n4948), .A2(n4938), .ZN(n4992) );
  CKND2D0 U4724 ( .A1(n4982), .A2(n5011), .ZN(n4938) );
  AO21D0 U4725 ( .A1(n4979), .A2(n5012), .B(n3527), .Z(n5011) );
  OA21D0 U4726 ( .A1(n5013), .A2(n5014), .B(n5015), .Z(n4982) );
  OAI211D0 U4727 ( .A1(n5016), .A2(n3527), .B(n4983), .C(n4976), .ZN(n4948) );
  OA211D0 U4728 ( .A1(n3578), .A2(n3527), .B(n3572), .C(n3569), .Z(n4976) );
  AN2D0 U4729 ( .A1(n5017), .A2(n5018), .Z(n3578) );
  AN2D0 U4730 ( .A1(n3262), .A2(n5019), .Z(n4983) );
  AN4D0 U4731 ( .A1(n3571), .A2(n5020), .A3(n3538), .A4(n5021), .Z(n3262) );
  NR2D0 U4732 ( .A1(n5022), .A2(n3545), .ZN(n5021) );
  CKND0 U4733 ( .I(n4978), .ZN(n5016) );
  ND4D0 U4734 ( .A1(n5023), .A2(n5024), .A3(n5025), .A4(n5026), .ZN(n4978) );
  CKND0 U4735 ( .I(n4774), .ZN(n4769) );
  OAI221D0 U4736 ( .A1(n5027), .A2(n5028), .B1(n5029), .B2(n3527), .C(n5030), 
        .ZN(n4774) );
  AOI221D0 U4737 ( .A1(n5031), .A2(n5032), .B1(n3550), .B2(n5033), .C(n5034), 
        .ZN(n5029) );
  OAI211D0 U4738 ( .A1(n5027), .A2(n5035), .B(n3581), .C(n5036), .ZN(n5033) );
  AOI21D0 U4739 ( .A1(n3531), .A2(n5037), .B(n3586), .ZN(n5036) );
  CKND0 U4740 ( .I(n5038), .ZN(n3586) );
  INR4D0 U4741 ( .A1(n5039), .B1(n5040), .B2(n4963), .B3(n5041), .ZN(n5035) );
  ND4D0 U4742 ( .A1(n3590), .A2(n5042), .A3(n3535), .A4(n3537), .ZN(n5040) );
  CKND0 U4743 ( .I(n4966), .ZN(n3590) );
  CKND2D0 U4744 ( .A1(n5043), .A2(n4970), .ZN(n5031) );
  INR2D0 U4745 ( .A1(n5044), .B1(n5045), .ZN(n4970) );
  INR3D0 U4746 ( .A1(n5046), .B1(n4953), .B2(n4971), .ZN(n5028) );
  ND3D0 U4747 ( .A1(n5047), .A2(n5020), .A3(n5048), .ZN(n4971) );
  CKND0 U4748 ( .I(n4797), .ZN(n4792) );
  OAI221D0 U4749 ( .A1(n5049), .A2(n5050), .B1(n5051), .B2(n3527), .C(n5052), 
        .ZN(n4797) );
  AOI221D0 U4750 ( .A1(n5053), .A2(n5054), .B1(n3550), .B2(n5055), .C(n5045), 
        .ZN(n5051) );
  CKND2D0 U4751 ( .A1(n3554), .A2(n3548), .ZN(n5045) );
  IND4D0 U4752 ( .A1(n3587), .B1(n5056), .B2(n5057), .B3(n3585), .ZN(n5055) );
  OAI31D0 U4753 ( .A1(n5058), .A2(n4968), .A3(n5059), .B(n5054), .ZN(n5057) );
  ND3D0 U4754 ( .A1(n5060), .A2(n5038), .A3(n3535), .ZN(n4968) );
  AN2D0 U4755 ( .A1(n3310), .A2(n5061), .Z(n3535) );
  ND3D0 U4756 ( .A1(n3537), .A2(n3581), .A3(n5062), .ZN(n5058) );
  OAI21D0 U4757 ( .A1(n5063), .A2(n4966), .B(n3531), .ZN(n5056) );
  IAO21D0 U4758 ( .A1(n4963), .A2(n4965), .B(n5049), .ZN(n5063) );
  ND3D0 U4759 ( .A1(n3591), .A2(n5064), .A3(n5042), .ZN(n4965) );
  CKND0 U4760 ( .I(n3532), .ZN(n5042) );
  ND4D0 U4761 ( .A1(n5065), .A2(n4988), .A3(n5066), .A4(n4987), .ZN(n3532) );
  CKND0 U4762 ( .I(n5067), .ZN(n4987) );
  NR2D0 U4763 ( .A1(n5068), .A2(n5069), .ZN(n5066) );
  ND3D0 U4764 ( .A1(n4969), .A2(n5044), .A3(n5043), .ZN(n5053) );
  CKND0 U4765 ( .I(n4957), .ZN(n5043) );
  CKND2D0 U4766 ( .A1(n3546), .A2(n3547), .ZN(n4957) );
  AN3D0 U4767 ( .A1(n5070), .A2(n5071), .A3(n3526), .Z(n5044) );
  AN3D0 U4768 ( .A1(n5072), .A2(n5073), .A3(n5074), .Z(n3526) );
  CKND0 U4769 ( .I(n5075), .ZN(n5072) );
  CKND0 U4770 ( .I(n5034), .ZN(n4969) );
  CKND2D0 U4771 ( .A1(n3597), .A2(n3598), .ZN(n5034) );
  NR2D0 U4772 ( .A1(n5076), .A2(n3530), .ZN(n5050) );
  CKND0 U4773 ( .I(n4830), .ZN(n4818) );
  OAI221D0 U4774 ( .A1(n5077), .A2(n5078), .B1(n5079), .B2(n3527), .C(n5080), 
        .ZN(n4830) );
  CKND0 U4775 ( .I(n3530), .ZN(n5080) );
  CKND2D0 U4776 ( .A1(n5020), .A2(n5081), .ZN(n3530) );
  ND4D0 U4777 ( .A1(n5082), .A2(n5083), .A3(n5084), .A4(n5085), .ZN(n5020) );
  CKND2D0 U4778 ( .A1(n5086), .A2(n5087), .ZN(n3527) );
  AOI221D0 U4779 ( .A1(n5088), .A2(n5089), .B1(n3550), .B2(n5090), .C(n5075), 
        .ZN(n5079) );
  CKND2D0 U4780 ( .A1(n5025), .A2(n5026), .ZN(n5075) );
  ND4D0 U4781 ( .A1(n5091), .A2(n5061), .A3(n5092), .A4(n3537), .ZN(n5090) );
  OAI21D0 U4782 ( .A1(n5069), .A2(n5068), .B(n3531), .ZN(n5092) );
  CKND0 U4783 ( .I(n3556), .ZN(n3531) );
  CKND2D0 U4784 ( .A1(n3559), .A2(n5093), .ZN(n3556) );
  CKND0 U4785 ( .I(n5094), .ZN(n5068) );
  CKND0 U4786 ( .I(n5095), .ZN(n5069) );
  OAI21D0 U4787 ( .A1(n5096), .A2(n5097), .B(n5089), .ZN(n5091) );
  IND4D0 U4788 ( .A1(n5041), .B1(n3555), .B2(n5039), .B3(n3591), .ZN(n5097) );
  CKND0 U4789 ( .I(n5037), .ZN(n3591) );
  CKND2D0 U4790 ( .A1(n5006), .A2(n5098), .ZN(n5037) );
  NR2D0 U4791 ( .A1(n5059), .A2(n3561), .ZN(n5039) );
  CKND0 U4792 ( .I(n3585), .ZN(n3561) );
  IND3D0 U4793 ( .A1(n3534), .B1(n5099), .B2(n4959), .ZN(n5059) );
  NR4D0 U4794 ( .A1(n4963), .A2(n4966), .A3(n3340), .A4(n5067), .ZN(n3555) );
  CKND2D0 U4795 ( .A1(n5005), .A2(n5100), .ZN(n4966) );
  CKND2D0 U4796 ( .A1(n5101), .A2(n5102), .ZN(n4963) );
  ND4D0 U4797 ( .A1(n3564), .A2(n5060), .A3(n5064), .A4(n4150), .ZN(n5041) );
  ND4D0 U4798 ( .A1(n5065), .A2(n3310), .A3(n3581), .A4(n5038), .ZN(n5096) );
  CKND0 U4799 ( .I(n3594), .ZN(n5065) );
  CKND2D0 U4800 ( .A1(n5103), .A2(n3339), .ZN(n3594) );
  CKND0 U4801 ( .I(n3576), .ZN(n3550) );
  ND3D0 U4802 ( .A1(n5104), .A2(n5105), .A3(n5106), .ZN(n3576) );
  AOI211D0 U4803 ( .A1(n5107), .A2(n5108), .B(n5109), .C(n5110), .ZN(n5106) );
  OAI22D0 U4804 ( .A1(n4302), .A2(n4940), .B1(n4043), .B2(n4999), .ZN(n5108)
         );
  IND3D0 U4805 ( .A1(n3266), .B1(n5023), .B2(n5073), .ZN(n5088) );
  INR2D0 U4806 ( .A1(n5052), .B1(n5076), .ZN(n5078) );
  OR2D0 U4807 ( .A1(n4972), .A2(n4953), .Z(n5076) );
  CKND2D0 U4808 ( .A1(n3538), .A2(n3539), .ZN(n4953) );
  IND3D0 U4809 ( .A1(n5111), .B1(n5112), .B2(n5113), .ZN(n3538) );
  CKND2D0 U4810 ( .A1(n5046), .A2(n5030), .ZN(n4972) );
  AN2D0 U4811 ( .A1(n3571), .A2(n3570), .Z(n5030) );
  OR2D0 U4812 ( .A1(n5112), .A2(n5022), .Z(n3571) );
  INR3D0 U4813 ( .A1(n5114), .B1(n5022), .B2(n3529), .ZN(n5046) );
  CKND2D0 U4814 ( .A1(n3260), .A2(n5115), .ZN(n3529) );
  AN3D0 U4815 ( .A1(n3572), .A2(n5015), .A3(n4996), .Z(n3260) );
  ND3D0 U4816 ( .A1(n5086), .A2(n5084), .A3(n5116), .ZN(n4996) );
  AOI211D0 U4817 ( .A1(n4934), .A2(n3946), .B(n4999), .C(n3373), .ZN(n5116) );
  ND4D0 U4818 ( .A1(n5086), .A2(n5084), .A3(n4934), .A4(n3946), .ZN(n5015) );
  OA211D0 U4819 ( .A1(n5117), .A2(n5118), .B(n5085), .C(n5083), .Z(n5086) );
  CKND0 U4820 ( .I(n5119), .ZN(n5085) );
  AOI21D0 U4821 ( .A1(n4974), .A2(n4014), .B(n5082), .ZN(n5117) );
  ND4D0 U4822 ( .A1(n5084), .A2(n4974), .A3(n5083), .A4(n5120), .ZN(n3572) );
  NR3D0 U4823 ( .A1(n3372), .A2(n5082), .A3(n5119), .ZN(n5120) );
  INR2D0 U4824 ( .A1(n4016), .B1(n5089), .ZN(n5082) );
  CKND0 U4825 ( .I(n5113), .ZN(n5022) );
  INR2D0 U4826 ( .A1(n3540), .B1(n3545), .ZN(n5052) );
  CKND0 U4827 ( .I(n5047), .ZN(n3545) );
  CKND2D0 U4828 ( .A1(n5119), .A2(n5083), .ZN(n5047) );
  AN3D0 U4829 ( .A1(n5111), .A2(n5113), .A3(n5112), .Z(n5083) );
  IND3D0 U4830 ( .A1(n3894), .B1(n5027), .B2(n5084), .ZN(n5112) );
  CKND2D0 U4831 ( .A1(n5084), .A2(n3893), .ZN(n5113) );
  ND3D0 U4832 ( .A1(n4949), .A2(n4019), .A3(n5084), .ZN(n5111) );
  CKND0 U4833 ( .I(n5118), .ZN(n5084) );
  NR3D0 U4834 ( .A1(n5054), .A2(n4011), .A3(n5118), .ZN(n5119) );
  CKND2D0 U4835 ( .A1(n3261), .A2(n5121), .ZN(n5118) );
  AN2D0 U4836 ( .A1(n5019), .A2(n5115), .Z(n3261) );
  OA211D0 U4837 ( .A1(n5013), .A2(n5014), .B(n4995), .C(n3569), .Z(n5115) );
  IND3D0 U4838 ( .A1(n5122), .B1(n5123), .B2(n5124), .ZN(n3569) );
  ND4D0 U4839 ( .A1(n5087), .A2(n5121), .A3(n5125), .A4(n4991), .ZN(n4995) );
  AN2D0 U4840 ( .A1(n5014), .A2(n4028), .Z(n5125) );
  CKND0 U4841 ( .I(n5013), .ZN(n5087) );
  ND3D0 U4842 ( .A1(n4934), .A2(n4034), .A3(n5121), .ZN(n5014) );
  ND3D0 U4843 ( .A1(n5122), .A2(n5123), .A3(n5124), .ZN(n5013) );
  ND3D0 U4844 ( .A1(n4974), .A2(n4029), .A3(n5121), .ZN(n5122) );
  AN4D0 U4845 ( .A1(n5048), .A2(n5114), .A3(n3539), .A4(n3570), .Z(n5019) );
  IND2D0 U4846 ( .A1(n5126), .B1(n5114), .ZN(n3570) );
  IND2D0 U4847 ( .A1(n5127), .B1(n5128), .ZN(n3539) );
  AN2D0 U4848 ( .A1(n5081), .A2(n3540), .Z(n5048) );
  IND2D0 U4849 ( .A1(n5123), .B1(n5124), .ZN(n5081) );
  AN3D0 U4850 ( .A1(n5127), .A2(n5129), .A3(n5128), .Z(n5124) );
  ND3D0 U4851 ( .A1(n5077), .A2(n4033), .A3(n5121), .ZN(n5123) );
  IND3D0 U4852 ( .A1(n5129), .B1(n5128), .B2(n5127), .ZN(n3540) );
  ND3D0 U4853 ( .A1(n4949), .A2(n4037), .A3(n5121), .ZN(n5127) );
  AN2D0 U4854 ( .A1(n5126), .A2(n5114), .Z(n5128) );
  CKND2D0 U4855 ( .A1(n5121), .A2(n4035), .ZN(n5114) );
  ND3D0 U4856 ( .A1(n5027), .A2(n4352), .A3(n5121), .ZN(n5126) );
  ND3D0 U4857 ( .A1(n5049), .A2(n4038), .A3(n5121), .ZN(n5129) );
  INR2D0 U4858 ( .A1(n5107), .B1(n3264), .ZN(n5121) );
  ND3D0 U4859 ( .A1(n5023), .A2(n5025), .A3(n5073), .ZN(n3264) );
  AN2D0 U4860 ( .A1(n4981), .A2(n5018), .Z(n5073) );
  IND3D0 U4861 ( .A1(n5130), .B1(n5131), .B2(n5132), .ZN(n5018) );
  AN2D0 U4862 ( .A1(n5012), .A2(n4997), .Z(n4981) );
  ND3D0 U4863 ( .A1(n5104), .A2(n5107), .A3(n5133), .ZN(n4997) );
  AOI211D0 U4864 ( .A1(n4934), .A2(n4042), .B(n4999), .C(n4043), .ZN(n5133) );
  ND4D0 U4865 ( .A1(n5104), .A2(n5107), .A3(n4934), .A4(n4042), .ZN(n5012) );
  AN3D0 U4866 ( .A1(n5130), .A2(n5132), .A3(n5131), .Z(n5104) );
  ND3D0 U4867 ( .A1(n4974), .A2(n4047), .A3(n5107), .ZN(n5130) );
  IND2D0 U4868 ( .A1(n5132), .B1(n5131), .ZN(n5025) );
  AN3D0 U4869 ( .A1(n5134), .A2(n5135), .A3(n5136), .Z(n5131) );
  ND3D0 U4870 ( .A1(n5077), .A2(n4053), .A3(n5107), .ZN(n5132) );
  AN4D0 U4871 ( .A1(n3554), .A2(n5070), .A3(n3546), .A4(n3597), .Z(n5023) );
  IND2D0 U4872 ( .A1(n5137), .B1(n5070), .ZN(n3597) );
  IND2D0 U4873 ( .A1(n5134), .B1(n5136), .ZN(n3546) );
  IND3D0 U4874 ( .A1(n5135), .B1(n5136), .B2(n5134), .ZN(n3554) );
  ND3D0 U4875 ( .A1(n4949), .A2(n4052), .A3(n5107), .ZN(n5134) );
  AN2D0 U4876 ( .A1(n5137), .A2(n5070), .Z(n5136) );
  CKND2D0 U4877 ( .A1(n5107), .A2(n4049), .ZN(n5070) );
  ND3D0 U4878 ( .A1(n5027), .A2(n4361), .A3(n5107), .ZN(n5137) );
  ND3D0 U4879 ( .A1(n5049), .A2(n4051), .A3(n5107), .ZN(n5135) );
  INR3D0 U4880 ( .A1(n5138), .B1(n3266), .B2(n3265), .ZN(n5107) );
  CKND0 U4881 ( .I(n5026), .ZN(n3265) );
  IND2D0 U4882 ( .A1(n5139), .B1(n5140), .ZN(n5026) );
  CKND2D0 U4883 ( .A1(n5024), .A2(n5074), .ZN(n3266) );
  AN3D0 U4884 ( .A1(n5017), .A2(n4980), .A3(n4979), .Z(n5074) );
  CKND2D0 U4885 ( .A1(n5109), .A2(n5105), .ZN(n4979) );
  CKND0 U4886 ( .I(n5141), .ZN(n5109) );
  ND3D0 U4887 ( .A1(n5110), .A2(n5141), .A3(n5105), .ZN(n4980) );
  AN3D0 U4888 ( .A1(n5142), .A2(n5139), .A3(n5140), .Z(n5105) );
  ND3D0 U4889 ( .A1(n4934), .A2(n4062), .A3(n5138), .ZN(n5141) );
  AN3D0 U4890 ( .A1(n4991), .A2(n4060), .A3(n5138), .Z(n5110) );
  IND3D0 U4891 ( .A1(n5142), .B1(n5140), .B2(n5139), .ZN(n5017) );
  ND3D0 U4892 ( .A1(n5077), .A2(n4066), .A3(n5138), .ZN(n5139) );
  AN3D0 U4893 ( .A1(n5143), .A2(n5144), .A3(n5145), .Z(n5140) );
  ND3D0 U4894 ( .A1(n4974), .A2(n4065), .A3(n5138), .ZN(n5142) );
  AN4D0 U4895 ( .A1(n3548), .A2(n5071), .A3(n3547), .A4(n3598), .Z(n5024) );
  IND2D0 U4896 ( .A1(n5146), .B1(n5071), .ZN(n3598) );
  IND2D0 U4897 ( .A1(n5143), .B1(n5145), .ZN(n3547) );
  IND3D0 U4898 ( .A1(n5144), .B1(n5145), .B2(n5143), .ZN(n3548) );
  ND3D0 U4899 ( .A1(n4949), .A2(n4069), .A3(n5138), .ZN(n5143) );
  AN2D0 U4900 ( .A1(n5146), .A2(n5071), .Z(n5145) );
  CKND2D0 U4901 ( .A1(n5138), .A2(n4067), .ZN(n5071) );
  ND3D0 U4902 ( .A1(n5027), .A2(n4371), .A3(n5138), .ZN(n5146) );
  ND3D0 U4903 ( .A1(n5049), .A2(n4070), .A3(n5138), .ZN(n5144) );
  AN2D0 U4904 ( .A1(n3341), .A2(n5147), .Z(n5138) );
  NR3D0 U4905 ( .A1(n3534), .A2(n3562), .A3(n4967), .ZN(n3341) );
  ND4D0 U4906 ( .A1(n3585), .A2(n5099), .A3(n3537), .A4(n3581), .ZN(n4967) );
  IND2D0 U4907 ( .A1(n5148), .B1(n5099), .ZN(n3581) );
  IND2D0 U4908 ( .A1(n5149), .B1(n5150), .ZN(n3537) );
  IND3D0 U4909 ( .A1(n5151), .B1(n5152), .B2(n5153), .ZN(n3585) );
  CKND0 U4910 ( .I(n4959), .ZN(n3562) );
  IND2D0 U4911 ( .A1(n5153), .B1(n5152), .ZN(n4959) );
  CKND2D0 U4912 ( .A1(n3557), .A2(n3582), .ZN(n3534) );
  IND3D0 U4913 ( .A1(n5154), .B1(n5150), .B2(n5149), .ZN(n3582) );
  AN2D0 U4914 ( .A1(n5008), .A2(n3584), .Z(n3557) );
  ND3D0 U4915 ( .A1(n3559), .A2(n5147), .A3(n5155), .ZN(n3584) );
  AOI211D0 U4916 ( .A1(n4934), .A2(n4076), .B(n4999), .C(n4077), .ZN(n5155) );
  ND4D0 U4917 ( .A1(n3559), .A2(n5147), .A3(n4934), .A4(n4076), .ZN(n5008) );
  CKND0 U4918 ( .I(n3536), .ZN(n3559) );
  ND3D0 U4919 ( .A1(n5154), .A2(n5149), .A3(n5150), .ZN(n3536) );
  AN3D0 U4920 ( .A1(n5151), .A2(n5153), .A3(n5152), .Z(n5150) );
  AN2D0 U4921 ( .A1(n5148), .A2(n5099), .Z(n5152) );
  CKND2D0 U4922 ( .A1(n5147), .A2(n4079), .ZN(n5099) );
  ND3D0 U4923 ( .A1(n5027), .A2(n5156), .A3(n5147), .ZN(n5148) );
  ND3D0 U4924 ( .A1(n4949), .A2(n4082), .A3(n5147), .ZN(n5153) );
  ND3D0 U4925 ( .A1(n5049), .A2(n4081), .A3(n5147), .ZN(n5151) );
  ND3D0 U4926 ( .A1(n5077), .A2(n4083), .A3(n5147), .ZN(n5149) );
  ND3D0 U4927 ( .A1(n4974), .A2(n5157), .A3(n5147), .ZN(n5154) );
  AN3D0 U4928 ( .A1(n5158), .A2(n3311), .A3(n3310), .Z(n5147) );
  NR2D0 U4929 ( .A1(n3563), .A2(n3588), .ZN(n3310) );
  CKND0 U4930 ( .I(n5003), .ZN(n3588) );
  IND3D0 U4931 ( .A1(n5159), .B1(n5160), .B2(n5161), .ZN(n5003) );
  CKND2D0 U4932 ( .A1(n5007), .A2(n3580), .ZN(n3563) );
  ND3D0 U4933 ( .A1(n5093), .A2(n5158), .A3(n5162), .ZN(n3580) );
  AOI211D0 U4934 ( .A1(n4934), .A2(n4097), .B(n4999), .C(n4092), .ZN(n5162) );
  ND4D0 U4935 ( .A1(n5093), .A2(n5158), .A3(n4934), .A4(n4097), .ZN(n5007) );
  CKND0 U4936 ( .I(n3593), .ZN(n5093) );
  ND3D0 U4937 ( .A1(n5159), .A2(n5161), .A3(n5160), .ZN(n3593) );
  ND3D0 U4938 ( .A1(n4974), .A2(n4087), .A3(n5158), .ZN(n5159) );
  AN4D0 U4939 ( .A1(n3564), .A2(n5060), .A3(n5061), .A4(n5038), .Z(n3311) );
  IND2D0 U4940 ( .A1(n5163), .B1(n5060), .ZN(n5038) );
  IND2D0 U4941 ( .A1(n5161), .B1(n5160), .ZN(n5061) );
  AN3D0 U4942 ( .A1(n5164), .A2(n5165), .A3(n5166), .Z(n5160) );
  ND3D0 U4943 ( .A1(n5077), .A2(n4096), .A3(n5158), .ZN(n5161) );
  NR2D0 U4944 ( .A1(n3587), .A2(n4962), .ZN(n3564) );
  CKND0 U4945 ( .I(n5062), .ZN(n4962) );
  CKND2D0 U4946 ( .A1(n5167), .A2(n5166), .ZN(n5062) );
  INR3D0 U4947 ( .A1(n5166), .B1(n5167), .B2(n5165), .ZN(n3587) );
  ND3D0 U4948 ( .A1(n5049), .A2(n4101), .A3(n5158), .ZN(n5165) );
  CKND0 U4949 ( .I(n5164), .ZN(n5167) );
  ND3D0 U4950 ( .A1(n4949), .A2(n4100), .A3(n5158), .ZN(n5164) );
  AN2D0 U4951 ( .A1(n5163), .A2(n5060), .Z(n5166) );
  CKND2D0 U4952 ( .A1(n5158), .A2(n4098), .ZN(n5060) );
  ND3D0 U4953 ( .A1(n5027), .A2(n5168), .A3(n5158), .ZN(n5163) );
  AN4D0 U4954 ( .A1(n3338), .A2(n4988), .A3(n5169), .A4(n3339), .Z(n5158) );
  ND3D0 U4955 ( .A1(n5170), .A2(n5169), .A3(n5171), .ZN(n3339) );
  AOI211D0 U4956 ( .A1(n5077), .A2(n4115), .B(n4985), .C(n4114), .ZN(n5171) );
  CKND0 U4957 ( .I(n3340), .ZN(n4988) );
  CKND2D0 U4958 ( .A1(n5010), .A2(n5002), .ZN(n3340) );
  ND3D0 U4959 ( .A1(n5172), .A2(n5169), .A3(n5173), .ZN(n5002) );
  AOI211D0 U4960 ( .A1(n4934), .A2(n4106), .B(n4999), .C(n4107), .ZN(n5173) );
  ND4D0 U4961 ( .A1(n5172), .A2(n5169), .A3(n4934), .A4(n4106), .ZN(n5010) );
  OA221D0 U4962 ( .A1(n4397), .A2(n5089), .B1(n4114), .B2(n4985), .C(n5170), 
        .Z(n5172) );
  AN4D0 U4963 ( .A1(n5098), .A2(n5064), .A3(n5095), .A4(n5174), .Z(n3338) );
  AN2D0 U4964 ( .A1(n5100), .A2(n5101), .Z(n5174) );
  IND2D0 U4965 ( .A1(n5175), .B1(n5176), .ZN(n5101) );
  IND3D0 U4966 ( .A1(n5177), .B1(n5176), .B2(n5175), .ZN(n5100) );
  ND4D0 U4967 ( .A1(n5170), .A2(n5169), .A3(n5077), .A4(n4115), .ZN(n5095) );
  AN3D0 U4968 ( .A1(n5175), .A2(n5177), .A3(n5176), .Z(n5170) );
  AN2D0 U4969 ( .A1(n5178), .A2(n5064), .Z(n5176) );
  ND3D0 U4970 ( .A1(n5049), .A2(n4104), .A3(n5169), .ZN(n5177) );
  ND3D0 U4971 ( .A1(n4949), .A2(n4113), .A3(n5169), .ZN(n5175) );
  CKND0 U4972 ( .I(n4955), .ZN(n4949) );
  IND2D0 U4973 ( .A1(n5178), .B1(n5064), .ZN(n5098) );
  CKND2D0 U4974 ( .A1(n5169), .A2(n4112), .ZN(n5064) );
  ND3D0 U4975 ( .A1(n5027), .A2(n4111), .A3(n5169), .ZN(n5178) );
  AN4D0 U4976 ( .A1(n5006), .A2(n5103), .A3(n5005), .A4(n5179), .Z(n5169) );
  NR2D0 U4977 ( .A1(n5067), .A2(n5004), .ZN(n5179) );
  ND3D0 U4978 ( .A1(n4150), .A2(n5102), .A3(n5094), .ZN(n5004) );
  IND3D0 U4979 ( .A1(n5180), .B1(n5181), .B2(n5182), .ZN(n5094) );
  CKND2D0 U4980 ( .A1(n5183), .A2(n4150), .ZN(n5102) );
  CKND2D0 U4981 ( .A1(n5001), .A2(n5009), .ZN(n5067) );
  ND3D0 U4982 ( .A1(n5184), .A2(n4121), .A3(n4934), .ZN(n5009) );
  ND4D0 U4983 ( .A1(n4991), .A2(n5184), .A3(n4119), .A4(n5185), .ZN(n5001) );
  CKND2D0 U4984 ( .A1(n4934), .A2(n4121), .ZN(n5185) );
  CKND0 U4985 ( .I(n4940), .ZN(n4934) );
  OAI221D0 U4986 ( .A1(n5186), .A2(n5187), .B1(n5188), .B2(n3442), .C(n5189), 
        .ZN(n4940) );
  CKND0 U4987 ( .I(n5190), .ZN(n5189) );
  AOI221D0 U4988 ( .A1(n5191), .A2(n5192), .B1(n5193), .B2(n5194), .C(n5195), 
        .ZN(n5188) );
  OAI211D0 U4989 ( .A1(n5186), .A2(n5196), .B(n5197), .C(n5198), .ZN(n5194) );
  CKND0 U4990 ( .I(n5199), .ZN(n5196) );
  CKND2D0 U4991 ( .A1(n5200), .A2(n5201), .ZN(n5191) );
  NR2D0 U4992 ( .A1(n5202), .A2(n5203), .ZN(n5187) );
  OA21D0 U4993 ( .A1(n4146), .A2(n4985), .B(n5204), .Z(n5184) );
  CKND0 U4994 ( .I(n4999), .ZN(n4991) );
  OAI221D0 U4995 ( .A1(n5205), .A2(n5206), .B1(n5201), .B2(n3442), .C(n5207), 
        .ZN(n4999) );
  CKND0 U4996 ( .I(n5202), .ZN(n5207) );
  OAI21D0 U4997 ( .A1(n3466), .A2(n5208), .B(n3455), .ZN(n5202) );
  AN2D0 U4998 ( .A1(n5209), .A2(n5210), .Z(n3466) );
  OA211D0 U4999 ( .A1(n5211), .A2(n3438), .B(n3474), .C(n3468), .Z(n5201) );
  NR2D0 U5000 ( .A1(n3483), .A2(n3485), .ZN(n5211) );
  CKND0 U5001 ( .I(n5212), .ZN(n3485) );
  CKND0 U5002 ( .I(n5213), .ZN(n3483) );
  AOI211D0 U5003 ( .A1(n5214), .A2(n5215), .B(n5190), .C(n5203), .ZN(n5206) );
  OAI211D0 U5004 ( .A1(n5216), .A2(n5208), .B(n5217), .C(n5218), .ZN(n5203) );
  CKND0 U5005 ( .I(n5219), .ZN(n5216) );
  CKND2D0 U5006 ( .A1(n5220), .A2(n5221), .ZN(n5190) );
  AO21D0 U5007 ( .A1(n5222), .A2(n5223), .B(n5208), .Z(n5221) );
  ND4D0 U5008 ( .A1(n5197), .A2(n5198), .A3(n5200), .A4(n5224), .ZN(n5215) );
  NR2D0 U5009 ( .A1(n5195), .A2(n5199), .ZN(n5224) );
  CKND2D0 U5010 ( .A1(n5225), .A2(n3480), .ZN(n5199) );
  CKND2D0 U5011 ( .A1(n5226), .A2(n5227), .ZN(n5195) );
  AN4D0 U5012 ( .A1(n5228), .A2(n5229), .A3(n5230), .A4(n3439), .Z(n5200) );
  CKND0 U5013 ( .I(n3442), .ZN(n5214) );
  CKND2D0 U5014 ( .A1(n5180), .A2(n5181), .ZN(n5005) );
  ND3D0 U5015 ( .A1(n4974), .A2(n4144), .A3(n5204), .ZN(n5103) );
  INR3D0 U5016 ( .A1(n5181), .B1(n5182), .B2(n5180), .ZN(n5204) );
  NR2D0 U5017 ( .A1(n5054), .A2(n4457), .ZN(n5180) );
  NR2D0 U5018 ( .A1(n5089), .A2(n4456), .ZN(n5182) );
  INR2D0 U5019 ( .A1(n4150), .B1(n5183), .ZN(n5181) );
  NR2D0 U5020 ( .A1(n4955), .A2(n5231), .ZN(n5183) );
  OAI221D0 U5021 ( .A1(n5232), .A2(n5233), .B1(n5234), .B2(n5208), .C(n5235), 
        .ZN(n4955) );
  CKND0 U5022 ( .I(n5236), .ZN(n5235) );
  AOI221D0 U5023 ( .A1(n5237), .A2(n5238), .B1(n5239), .B2(n5240), .C(n5241), 
        .ZN(n5234) );
  OAI211D0 U5024 ( .A1(n5232), .A2(n5242), .B(n3439), .C(n5243), .ZN(n5240) );
  AOI21D0 U5025 ( .A1(n5193), .A2(n5244), .B(n5245), .ZN(n5243) );
  CKND0 U5026 ( .I(n5246), .ZN(n5245) );
  CKND2D0 U5027 ( .A1(n5247), .A2(n5248), .ZN(n5244) );
  OAI21D0 U5028 ( .A1(n5249), .A2(n3486), .B(n5238), .ZN(n5248) );
  INR4D0 U5029 ( .A1(n3454), .B1(n3477), .B2(n5250), .B3(n5251), .ZN(n5242) );
  CKND0 U5030 ( .I(n5252), .ZN(n3477) );
  IND2D0 U5031 ( .A1(n5253), .B1(n5254), .ZN(n5237) );
  NR2D0 U5032 ( .A1(n5255), .A2(n5256), .ZN(n5233) );
  IND2D0 U5033 ( .A1(n3937), .B1(n5027), .ZN(n5006) );
  CKND0 U5034 ( .I(n5032), .ZN(n5027) );
  OAI221D0 U5035 ( .A1(n5257), .A2(n5258), .B1(n5259), .B2(n5208), .C(n5260), 
        .ZN(n5032) );
  AOI221D0 U5036 ( .A1(n5261), .A2(n5262), .B1(n5239), .B2(n5263), .C(n5264), 
        .ZN(n5259) );
  OAI221D0 U5037 ( .A1(n5257), .A2(n5265), .B1(n3473), .B2(n5266), .C(n3469), 
        .ZN(n5263) );
  OAI33D0 U5038 ( .A1(n5262), .A2(n3484), .A3(n3475), .B1(n5267), .B2(n3486), 
        .B3(n5268), .ZN(n5266) );
  CKND2D0 U5039 ( .A1(n5269), .A2(n3315), .ZN(n5267) );
  NR2D0 U5040 ( .A1(n3452), .A2(n5270), .ZN(n5265) );
  CKND0 U5041 ( .I(n5271), .ZN(n3452) );
  IND3D0 U5042 ( .A1(n3447), .B1(n5272), .B2(n3431), .ZN(n5261) );
  INR3D0 U5043 ( .A1(n5273), .B1(n5236), .B2(n5255), .ZN(n5258) );
  ND3D0 U5044 ( .A1(n5274), .A2(n5275), .A3(n5276), .ZN(n5255) );
  CKND0 U5045 ( .I(n4985), .ZN(n4974) );
  OAI221D0 U5046 ( .A1(n5277), .A2(n3442), .B1(n5278), .B2(n5279), .C(n5218), 
        .ZN(n4985) );
  OA211D0 U5047 ( .A1(n3467), .A2(n5208), .B(n3462), .C(n3459), .Z(n5218) );
  AN2D0 U5048 ( .A1(n5280), .A2(n5281), .Z(n3467) );
  NR4D0 U5049 ( .A1(n5282), .A2(n3426), .A3(n3432), .A4(n5219), .ZN(n5279) );
  IND3D0 U5050 ( .A1(n3280), .B1(n5283), .B2(n5284), .ZN(n5219) );
  ND3D0 U5051 ( .A1(n5222), .A2(n5209), .A3(n5285), .ZN(n3432) );
  CKND2D0 U5052 ( .A1(n3455), .A2(n5220), .ZN(n3426) );
  OA21D0 U5053 ( .A1(n5286), .A2(n5287), .B(n5288), .Z(n5220) );
  AN2D0 U5054 ( .A1(n5289), .A2(n5290), .Z(n3455) );
  IND4D0 U5055 ( .A1(n3436), .B1(n5217), .B2(n5229), .B3(n3439), .ZN(n5282) );
  AN2D0 U5056 ( .A1(n3276), .A2(n5291), .Z(n5217) );
  AN4D0 U5057 ( .A1(n3461), .A2(n5275), .A3(n3420), .A4(n5292), .Z(n3276) );
  NR2D0 U5058 ( .A1(n5293), .A2(n3427), .ZN(n5292) );
  CKND2D0 U5059 ( .A1(n3424), .A2(n5239), .ZN(n3442) );
  CKND0 U5060 ( .I(n5208), .ZN(n3424) );
  AOI211D0 U5061 ( .A1(n5294), .A2(n5295), .B(n5296), .C(n5297), .ZN(n5277) );
  CKND0 U5062 ( .I(n5228), .ZN(n5296) );
  NR2D0 U5063 ( .A1(n3471), .A2(n3476), .ZN(n5228) );
  CKND0 U5064 ( .I(n5298), .ZN(n3476) );
  ND4D0 U5065 ( .A1(n5225), .A2(n5299), .A3(n5300), .A4(n5230), .ZN(n5294) );
  AN2D0 U5066 ( .A1(n5301), .A2(n5302), .Z(n5225) );
  CKND0 U5067 ( .I(n5054), .ZN(n5049) );
  OAI221D0 U5068 ( .A1(n5303), .A2(n5304), .B1(n5305), .B2(n5208), .C(n5306), 
        .ZN(n5054) );
  AOI221D0 U5069 ( .A1(n5307), .A2(n5308), .B1(n5239), .B2(n5309), .C(n5253), 
        .ZN(n5305) );
  CKND2D0 U5070 ( .A1(n3487), .A2(n3488), .ZN(n5253) );
  ND4D0 U5071 ( .A1(n5310), .A2(n5252), .A3(n5311), .A4(n3440), .ZN(n5309) );
  OAI31D0 U5072 ( .A1(n5312), .A2(n5251), .A3(n5313), .B(n5308), .ZN(n5311) );
  IND2D0 U5073 ( .A1(n3450), .B1(n5314), .ZN(n5251) );
  ND3D0 U5074 ( .A1(n5298), .A2(n5315), .A3(n5300), .ZN(n3450) );
  ND3D0 U5075 ( .A1(n5271), .A2(n3469), .A3(n5246), .ZN(n5312) );
  OAI21D0 U5076 ( .A1(n5316), .A2(n3486), .B(n5193), .ZN(n5310) );
  CKND0 U5077 ( .I(n3438), .ZN(n5193) );
  CKND2D0 U5078 ( .A1(n3433), .A2(n5317), .ZN(n3438) );
  AOI21D0 U5079 ( .A1(n5247), .A2(n5269), .B(n5303), .ZN(n5316) );
  CKND0 U5080 ( .I(n5249), .ZN(n5269) );
  CKND2D0 U5081 ( .A1(n3453), .A2(n5318), .ZN(n5249) );
  AN4D0 U5082 ( .A1(n5299), .A2(n3480), .A3(n5319), .A4(n5320), .Z(n3453) );
  CKND0 U5083 ( .I(n5268), .ZN(n5247) );
  IND2D0 U5084 ( .A1(n5241), .B1(n5254), .ZN(n5307) );
  INR2D0 U5085 ( .A1(n5321), .B1(n3447), .ZN(n5254) );
  CKND2D0 U5086 ( .A1(n5322), .A2(n5323), .ZN(n5241) );
  NR2D0 U5087 ( .A1(n5324), .A2(n3446), .ZN(n5304) );
  CKND0 U5088 ( .I(n5089), .ZN(n5077) );
  OAI221D0 U5089 ( .A1(n5325), .A2(n5326), .B1(n5327), .B2(n5208), .C(n5328), 
        .ZN(n5089) );
  CKND0 U5090 ( .I(n3446), .ZN(n5328) );
  CKND2D0 U5091 ( .A1(n5275), .A2(n5329), .ZN(n3446) );
  ND4D0 U5092 ( .A1(n5330), .A2(n5331), .A3(n5332), .A4(n5333), .ZN(n5275) );
  CKND2D0 U5093 ( .A1(n5334), .A2(n5335), .ZN(n5208) );
  AOI221D0 U5094 ( .A1(n5336), .A2(n5337), .B1(n5239), .B2(n5338), .C(n3447), 
        .ZN(n5327) );
  CKND2D0 U5095 ( .A1(n5339), .A2(n5340), .ZN(n3447) );
  OAI211D0 U5096 ( .A1(n5325), .A2(n5341), .B(n5319), .C(n5342), .ZN(n5338) );
  AN3D0 U5097 ( .A1(n5320), .A2(n5315), .A3(n5271), .Z(n5342) );
  NR4D0 U5098 ( .A1(n5343), .A2(n5344), .A3(n3434), .A4(n5270), .ZN(n5341) );
  IND2D0 U5099 ( .A1(n5313), .B1(n3440), .ZN(n5270) );
  ND3D0 U5100 ( .A1(n3439), .A2(n5345), .A3(n3454), .ZN(n5313) );
  ND3D0 U5101 ( .A1(n5246), .A2(n5252), .A3(n5300), .ZN(n3434) );
  CKND2D0 U5102 ( .A1(n3437), .A2(n5318), .ZN(n5344) );
  INR3D0 U5103 ( .A1(n4150), .B1(n3484), .B2(n5346), .ZN(n5318) );
  INR3D0 U5104 ( .A1(n5299), .B1(n3486), .B2(n5268), .ZN(n3437) );
  CKND2D0 U5105 ( .A1(n5347), .A2(n5348), .ZN(n5268) );
  CKND2D0 U5106 ( .A1(n5349), .A2(n5350), .ZN(n3486) );
  AN4D0 U5107 ( .A1(n5213), .A2(n5197), .A3(n5212), .A4(n5198), .Z(n5299) );
  ND4D0 U5108 ( .A1(n5314), .A2(n3480), .A3(n5298), .A4(n3469), .ZN(n5343) );
  CKND0 U5109 ( .I(n5297), .ZN(n3480) );
  CKND2D0 U5110 ( .A1(n5351), .A2(n5352), .ZN(n5297) );
  CKND0 U5111 ( .I(n3429), .ZN(n5239) );
  ND3D0 U5112 ( .A1(n5353), .A2(n5354), .A3(n5355), .ZN(n3429) );
  AOI211D0 U5113 ( .A1(n5356), .A2(n5357), .B(n5358), .C(n5359), .ZN(n5355) );
  OAI22D0 U5114 ( .A1(n4302), .A2(n5192), .B1(n4043), .B2(n5360), .ZN(n5357)
         );
  CKND2D0 U5115 ( .A1(n3431), .A2(n5321), .ZN(n5336) );
  INR2D0 U5116 ( .A1(n5272), .B1(n5264), .ZN(n5321) );
  CKND2D0 U5117 ( .A1(n3489), .A2(n3490), .ZN(n5264) );
  NR3D0 U5118 ( .A1(n3279), .A2(n5361), .A3(n3449), .ZN(n5272) );
  NR3D0 U5119 ( .A1(n5362), .A2(n5363), .A3(n5364), .ZN(n3431) );
  CKND0 U5120 ( .I(n5322), .ZN(n5363) );
  INR2D0 U5121 ( .A1(n5306), .B1(n5324), .ZN(n5326) );
  OR2D0 U5122 ( .A1(n5256), .A2(n5236), .Z(n5324) );
  CKND2D0 U5123 ( .A1(n3420), .A2(n3421), .ZN(n5236) );
  IND3D0 U5124 ( .A1(n5365), .B1(n5366), .B2(n5367), .ZN(n3420) );
  CKND2D0 U5125 ( .A1(n5273), .A2(n5260), .ZN(n5256) );
  AN2D0 U5126 ( .A1(n3461), .A2(n3460), .Z(n5260) );
  OR2D0 U5127 ( .A1(n5366), .A2(n5293), .Z(n3461) );
  INR3D0 U5128 ( .A1(n5368), .B1(n5293), .B2(n3445), .ZN(n5273) );
  CKND2D0 U5129 ( .A1(n3274), .A2(n5369), .ZN(n3445) );
  AN3D0 U5130 ( .A1(n3462), .A2(n5288), .A3(n5290), .Z(n3274) );
  ND3D0 U5131 ( .A1(n5334), .A2(n5332), .A3(n5370), .ZN(n5290) );
  AOI211D0 U5132 ( .A1(n5186), .A2(n3946), .B(n5360), .C(n3373), .ZN(n5370) );
  ND4D0 U5133 ( .A1(n5334), .A2(n5332), .A3(n5186), .A4(n3946), .ZN(n5288) );
  CKND0 U5134 ( .I(n3371), .ZN(n3946) );
  OA211D0 U5135 ( .A1(n5371), .A2(n5372), .B(n5333), .C(n5331), .Z(n5334) );
  CKND0 U5136 ( .I(n5373), .ZN(n5333) );
  AOI21D0 U5137 ( .A1(n5278), .A2(n4014), .B(n5330), .ZN(n5371) );
  ND4D0 U5138 ( .A1(n5332), .A2(n5278), .A3(n5331), .A4(n5374), .ZN(n3462) );
  NR3D0 U5139 ( .A1(n3372), .A2(n5330), .A3(n5373), .ZN(n5374) );
  INR2D0 U5140 ( .A1(n4016), .B1(n5337), .ZN(n5330) );
  CKND0 U5141 ( .I(n5367), .ZN(n5293) );
  INR2D0 U5142 ( .A1(n3422), .B1(n3427), .ZN(n5306) );
  CKND0 U5143 ( .I(n5274), .ZN(n3427) );
  CKND2D0 U5144 ( .A1(n5373), .A2(n5331), .ZN(n5274) );
  AN3D0 U5145 ( .A1(n5365), .A2(n5367), .A3(n5366), .Z(n5331) );
  IND3D0 U5146 ( .A1(n3894), .B1(n5257), .B2(n5332), .ZN(n5366) );
  CKND2D0 U5147 ( .A1(n5332), .A2(n3893), .ZN(n5367) );
  ND3D0 U5148 ( .A1(n5232), .A2(n4019), .A3(n5332), .ZN(n5365) );
  CKND0 U5149 ( .I(n5372), .ZN(n5332) );
  NR3D0 U5150 ( .A1(n5308), .A2(n4011), .A3(n5372), .ZN(n5373) );
  CKND2D0 U5151 ( .A1(n3275), .A2(n5375), .ZN(n5372) );
  AN2D0 U5152 ( .A1(n5291), .A2(n5369), .Z(n3275) );
  OA211D0 U5153 ( .A1(n5286), .A2(n5287), .B(n5289), .C(n3459), .Z(n5369) );
  IND3D0 U5154 ( .A1(n5376), .B1(n5377), .B2(n5378), .ZN(n3459) );
  ND4D0 U5155 ( .A1(n5335), .A2(n5375), .A3(n5379), .A4(n5205), .ZN(n5289) );
  AN2D0 U5156 ( .A1(n5287), .A2(n4028), .Z(n5379) );
  CKND0 U5157 ( .I(n5286), .ZN(n5335) );
  ND3D0 U5158 ( .A1(n5186), .A2(n4034), .A3(n5375), .ZN(n5287) );
  ND3D0 U5159 ( .A1(n5376), .A2(n5377), .A3(n5378), .ZN(n5286) );
  ND3D0 U5160 ( .A1(n5278), .A2(n4029), .A3(n5375), .ZN(n5376) );
  AN4D0 U5161 ( .A1(n5276), .A2(n5368), .A3(n3421), .A4(n3460), .Z(n5291) );
  IND2D0 U5162 ( .A1(n5380), .B1(n5368), .ZN(n3460) );
  IND2D0 U5163 ( .A1(n5381), .B1(n5382), .ZN(n3421) );
  AN2D0 U5164 ( .A1(n5329), .A2(n3422), .Z(n5276) );
  IND2D0 U5165 ( .A1(n5377), .B1(n5378), .ZN(n5329) );
  AN3D0 U5166 ( .A1(n5381), .A2(n5383), .A3(n5382), .Z(n5378) );
  ND3D0 U5167 ( .A1(n5325), .A2(n4033), .A3(n5375), .ZN(n5377) );
  IND3D0 U5168 ( .A1(n5383), .B1(n5382), .B2(n5381), .ZN(n3422) );
  ND3D0 U5169 ( .A1(n5232), .A2(n4037), .A3(n5375), .ZN(n5381) );
  AN2D0 U5170 ( .A1(n5380), .A2(n5368), .Z(n5382) );
  CKND2D0 U5171 ( .A1(n4035), .A2(n5375), .ZN(n5368) );
  ND3D0 U5172 ( .A1(n5257), .A2(n4352), .A3(n5375), .ZN(n5380) );
  ND3D0 U5173 ( .A1(n5303), .A2(n4038), .A3(n5375), .ZN(n5383) );
  INR2D0 U5174 ( .A1(n5356), .B1(n3278), .ZN(n5375) );
  CKND0 U5175 ( .I(n3351), .ZN(n3278) );
  INR2D0 U5176 ( .A1(n5284), .B1(n3449), .ZN(n3351) );
  CKND2D0 U5177 ( .A1(n5285), .A2(n5281), .ZN(n3449) );
  IND3D0 U5178 ( .A1(n5384), .B1(n5385), .B2(n5386), .ZN(n5281) );
  AN2D0 U5179 ( .A1(n5223), .A2(n5210), .Z(n5285) );
  ND3D0 U5180 ( .A1(n5353), .A2(n5356), .A3(n5387), .ZN(n5210) );
  AOI211D0 U5181 ( .A1(n5186), .A2(n4042), .B(n5360), .C(n4043), .ZN(n5387) );
  ND4D0 U5182 ( .A1(n5353), .A2(n5356), .A3(n5186), .A4(n4042), .ZN(n5223) );
  CKND0 U5183 ( .I(n4302), .ZN(n4042) );
  AN3D0 U5184 ( .A1(n5384), .A2(n5386), .A3(n5385), .Z(n5353) );
  ND3D0 U5185 ( .A1(n5278), .A2(n4047), .A3(n5356), .ZN(n5384) );
  CKND0 U5186 ( .I(n4045), .ZN(n4047) );
  AN4D0 U5187 ( .A1(n5339), .A2(n3489), .A3(n5322), .A4(n5388), .Z(n5284) );
  NR2D0 U5188 ( .A1(n5361), .A2(n5364), .ZN(n5388) );
  CKND0 U5189 ( .I(n3487), .ZN(n5364) );
  IND3D0 U5190 ( .A1(n5389), .B1(n5390), .B2(n5391), .ZN(n3487) );
  IND2D0 U5191 ( .A1(n5391), .B1(n5390), .ZN(n5322) );
  CKND2D0 U5192 ( .A1(n5392), .A2(n5393), .ZN(n3489) );
  IND2D0 U5193 ( .A1(n5386), .B1(n5385), .ZN(n5339) );
  AN3D0 U5194 ( .A1(n5391), .A2(n5389), .A3(n5390), .Z(n5385) );
  NR2D0 U5195 ( .A1(n5392), .A2(n5361), .ZN(n5390) );
  CKND0 U5196 ( .I(n5393), .ZN(n5361) );
  CKND2D0 U5197 ( .A1(n4049), .A2(n5356), .ZN(n5393) );
  AN3D0 U5198 ( .A1(n5356), .A2(n5257), .A3(n4361), .Z(n5392) );
  CKND0 U5199 ( .I(n4050), .ZN(n4361) );
  ND3D0 U5200 ( .A1(n5303), .A2(n4051), .A3(n5356), .ZN(n5389) );
  ND3D0 U5201 ( .A1(n5232), .A2(n4052), .A3(n5356), .ZN(n5391) );
  ND3D0 U5202 ( .A1(n5325), .A2(n4053), .A3(n5356), .ZN(n5386) );
  INR3D0 U5203 ( .A1(n5394), .B1(n3279), .B2(n3280), .ZN(n5356) );
  IND3D0 U5204 ( .A1(n5362), .B1(n5340), .B2(n3490), .ZN(n3280) );
  IND2D0 U5205 ( .A1(n5395), .B1(n5283), .ZN(n3490) );
  IND2D0 U5206 ( .A1(n5396), .B1(n5397), .ZN(n5340) );
  CKND2D0 U5207 ( .A1(n3488), .A2(n5323), .ZN(n5362) );
  IND2D0 U5208 ( .A1(n5398), .B1(n5399), .ZN(n5323) );
  IND3D0 U5209 ( .A1(n5400), .B1(n5399), .B2(n5398), .ZN(n3488) );
  IND2D0 U5210 ( .A1(n3448), .B1(n5283), .ZN(n3279) );
  ND3D0 U5211 ( .A1(n5280), .A2(n5209), .A3(n5222), .ZN(n3448) );
  CKND2D0 U5212 ( .A1(n5358), .A2(n5354), .ZN(n5222) );
  CKND0 U5213 ( .I(n5401), .ZN(n5358) );
  ND3D0 U5214 ( .A1(n5359), .A2(n5401), .A3(n5354), .ZN(n5209) );
  AN3D0 U5215 ( .A1(n5402), .A2(n5396), .A3(n5397), .Z(n5354) );
  ND3D0 U5216 ( .A1(n5186), .A2(n4062), .A3(n5394), .ZN(n5401) );
  AN3D0 U5217 ( .A1(n5205), .A2(n4060), .A3(n5394), .Z(n5359) );
  IND3D0 U5218 ( .A1(n5402), .B1(n5397), .B2(n5396), .ZN(n5280) );
  ND3D0 U5219 ( .A1(n5325), .A2(n4066), .A3(n5394), .ZN(n5396) );
  AN3D0 U5220 ( .A1(n5398), .A2(n5400), .A3(n5399), .Z(n5397) );
  AN2D0 U5221 ( .A1(n5395), .A2(n5283), .Z(n5399) );
  CKND2D0 U5222 ( .A1(n4067), .A2(n5394), .ZN(n5283) );
  ND3D0 U5223 ( .A1(n5257), .A2(n4371), .A3(n5394), .ZN(n5395) );
  CKND0 U5224 ( .I(n4068), .ZN(n4371) );
  ND3D0 U5225 ( .A1(n5303), .A2(n4070), .A3(n5394), .ZN(n5400) );
  ND3D0 U5226 ( .A1(n5232), .A2(n4069), .A3(n5394), .ZN(n5398) );
  ND3D0 U5227 ( .A1(n5278), .A2(n4065), .A3(n5394), .ZN(n5402) );
  AN2D0 U5228 ( .A1(n3353), .A2(n5403), .Z(n5394) );
  AN3D0 U5229 ( .A1(n3454), .A2(n3439), .A3(n5229), .Z(n3353) );
  CKND0 U5230 ( .I(n5250), .ZN(n5229) );
  ND4D0 U5231 ( .A1(n3440), .A2(n5345), .A3(n5271), .A4(n3469), .ZN(n5250) );
  IND2D0 U5232 ( .A1(n5404), .B1(n5345), .ZN(n3469) );
  CKND2D0 U5233 ( .A1(n5405), .A2(n5406), .ZN(n5271) );
  IND3D0 U5234 ( .A1(n5407), .B1(n5408), .B2(n5409), .ZN(n3440) );
  IND2D0 U5235 ( .A1(n5409), .B1(n5408), .ZN(n3439) );
  NR2D0 U5236 ( .A1(n3436), .A2(n3471), .ZN(n3454) );
  INR3D0 U5237 ( .A1(n5405), .B1(n5406), .B2(n5410), .ZN(n3471) );
  CKND0 U5238 ( .I(n5411), .ZN(n5406) );
  CKND2D0 U5239 ( .A1(n5227), .A2(n3474), .ZN(n3436) );
  ND3D0 U5240 ( .A1(n3433), .A2(n5403), .A3(n5412), .ZN(n3474) );
  AOI211D0 U5241 ( .A1(n5186), .A2(n4076), .B(n5360), .C(n4077), .ZN(n5412) );
  ND4D0 U5242 ( .A1(n3433), .A2(n5403), .A3(n5186), .A4(n4076), .ZN(n5227) );
  CKND0 U5243 ( .I(n3473), .ZN(n3433) );
  ND3D0 U5244 ( .A1(n5410), .A2(n5411), .A3(n5405), .ZN(n3473) );
  AN3D0 U5245 ( .A1(n5407), .A2(n5409), .A3(n5408), .Z(n5405) );
  AN2D0 U5246 ( .A1(n5404), .A2(n5345), .Z(n5408) );
  CKND2D0 U5247 ( .A1(n4079), .A2(n5403), .ZN(n5345) );
  ND3D0 U5248 ( .A1(n5257), .A2(n5156), .A3(n5403), .ZN(n5404) );
  CKND0 U5249 ( .I(n4080), .ZN(n5156) );
  ND3D0 U5250 ( .A1(n5232), .A2(n4082), .A3(n5403), .ZN(n5409) );
  ND3D0 U5251 ( .A1(n5303), .A2(n4081), .A3(n5403), .ZN(n5407) );
  CKND0 U5252 ( .I(n4004), .ZN(n4081) );
  ND3D0 U5253 ( .A1(n5325), .A2(n4083), .A3(n5403), .ZN(n5411) );
  ND3D0 U5254 ( .A1(n5278), .A2(n5157), .A3(n5403), .ZN(n5410) );
  AN2D0 U5255 ( .A1(n3315), .A2(n5413), .Z(n5403) );
  AN3D0 U5256 ( .A1(n5230), .A2(n5298), .A3(n5300), .Z(n3315) );
  AN2D0 U5257 ( .A1(n5226), .A2(n3468), .Z(n5300) );
  ND3D0 U5258 ( .A1(n5317), .A2(n5413), .A3(n5414), .ZN(n3468) );
  AOI211D0 U5259 ( .A1(n5186), .A2(n4097), .B(n5360), .C(n4092), .ZN(n5414) );
  ND4D0 U5260 ( .A1(n5317), .A2(n5413), .A3(n5186), .A4(n4097), .ZN(n5226) );
  CKND0 U5261 ( .I(n3482), .ZN(n5317) );
  ND3D0 U5262 ( .A1(n5415), .A2(n5416), .A3(n5417), .ZN(n3482) );
  IND3D0 U5263 ( .A1(n5416), .B1(n5417), .B2(n5415), .ZN(n5298) );
  ND3D0 U5264 ( .A1(n5278), .A2(n4087), .A3(n5413), .ZN(n5416) );
  AN4D0 U5265 ( .A1(n5314), .A2(n5246), .A3(n5252), .A4(n5315), .Z(n5230) );
  IND2D0 U5266 ( .A1(n5415), .B1(n5417), .ZN(n5315) );
  AN3D0 U5267 ( .A1(n5418), .A2(n5419), .A3(n5420), .Z(n5417) );
  ND3D0 U5268 ( .A1(n5325), .A2(n4096), .A3(n5413), .ZN(n5415) );
  IND3D0 U5269 ( .A1(n5419), .B1(n5420), .B2(n5418), .ZN(n5252) );
  ND3D0 U5270 ( .A1(n5303), .A2(n4101), .A3(n5413), .ZN(n5419) );
  IND2D0 U5271 ( .A1(n5418), .B1(n5420), .ZN(n5246) );
  AN2D0 U5272 ( .A1(n5421), .A2(n5422), .Z(n5420) );
  ND3D0 U5273 ( .A1(n5232), .A2(n4100), .A3(n5413), .ZN(n5418) );
  INR2D0 U5274 ( .A1(n5422), .B1(n3475), .ZN(n5314) );
  INR2D0 U5275 ( .A1(n5422), .B1(n5421), .ZN(n3475) );
  ND3D0 U5276 ( .A1(n5257), .A2(n5168), .A3(n5413), .ZN(n5421) );
  CKND0 U5277 ( .I(n4099), .ZN(n5168) );
  CKND2D0 U5278 ( .A1(n4098), .A2(n5413), .ZN(n5422) );
  AN2D0 U5279 ( .A1(n3352), .A2(n5423), .Z(n5413) );
  AN4D0 U5280 ( .A1(n5301), .A2(n5213), .A3(n5197), .A4(n5351), .Z(n3352) );
  ND3D0 U5281 ( .A1(n5278), .A2(n5424), .A3(n5425), .ZN(n5351) );
  ND3D0 U5282 ( .A1(n5186), .A2(n4106), .A3(n5426), .ZN(n5197) );
  ND4D0 U5283 ( .A1(n5426), .A2(n5205), .A3(n5427), .A4(n5428), .ZN(n5213) );
  CKND2D0 U5284 ( .A1(n5186), .A2(n4106), .ZN(n5428) );
  CKND0 U5285 ( .I(n5192), .ZN(n5186) );
  CKND0 U5286 ( .I(n5360), .ZN(n5205) );
  OA21D0 U5287 ( .A1(n4114), .A2(n5295), .B(n5425), .Z(n5426) );
  AN3D0 U5288 ( .A1(n5423), .A2(n5429), .A3(n5430), .Z(n5425) );
  AN4D0 U5289 ( .A1(n5347), .A2(n5350), .A3(n5431), .A4(n5319), .Z(n5301) );
  IND2D0 U5290 ( .A1(n5429), .B1(n5430), .ZN(n5319) );
  AN3D0 U5291 ( .A1(n5432), .A2(n5433), .A3(n5434), .Z(n5430) );
  ND3D0 U5292 ( .A1(n5325), .A2(n4115), .A3(n5423), .ZN(n5429) );
  NR2D0 U5293 ( .A1(n5346), .A2(n3484), .ZN(n5431) );
  NR2D0 U5294 ( .A1(n5435), .A2(n5346), .ZN(n3484) );
  IND3D0 U5295 ( .A1(n5433), .B1(n5434), .B2(n5432), .ZN(n5350) );
  ND3D0 U5296 ( .A1(n5303), .A2(n4104), .A3(n5423), .ZN(n5433) );
  CKND0 U5297 ( .I(n4110), .ZN(n4104) );
  IND2D0 U5298 ( .A1(n5432), .B1(n5434), .ZN(n5347) );
  INR2D0 U5299 ( .A1(n5435), .B1(n5346), .ZN(n5434) );
  AN2D0 U5300 ( .A1(n4112), .A2(n5423), .Z(n5346) );
  ND3D0 U5301 ( .A1(n4111), .A2(n5423), .A3(n5257), .ZN(n5435) );
  CKND0 U5302 ( .I(n5262), .ZN(n5257) );
  OAI211D0 U5303 ( .A1(n5436), .A2(n3318), .B(n3400), .C(n5437), .ZN(n5262) );
  NR2D0 U5304 ( .A1(n3396), .A2(n3414), .ZN(n5437) );
  OAI31D0 U5305 ( .A1(n5438), .A2(n4112), .A3(n5439), .B(n3937), .ZN(n3414) );
  IND2D0 U5306 ( .A1(n4149), .B1(n4150), .ZN(n3937) );
  OAI32D0 U5307 ( .A1(n4036), .A2(n4035), .A3(n5440), .B1(n3893), .B2(n5441), 
        .ZN(n3396) );
  CKND0 U5308 ( .I(n4283), .ZN(n3893) );
  CKND2D0 U5309 ( .A1(n5442), .A2(n5443), .ZN(n3400) );
  OAI33D0 U5310 ( .A1(n4068), .A2(n4067), .A3(n5444), .B1(n4050), .B2(n4049), 
        .B3(n5445), .ZN(n5443) );
  CKND0 U5311 ( .I(n3910), .ZN(n4049) );
  CKND0 U5312 ( .I(n3916), .ZN(n4067) );
  CKND0 U5313 ( .I(n3408), .ZN(n5436) );
  OAI33D0 U5314 ( .A1(n4099), .A2(n4098), .A3(n5446), .B1(n4080), .B2(n4079), 
        .B3(n5447), .ZN(n3408) );
  CKND0 U5315 ( .I(n3922), .ZN(n4079) );
  ND3D0 U5316 ( .A1(n5232), .A2(n4113), .A3(n5423), .ZN(n5432) );
  AN4D0 U5317 ( .A1(n5302), .A2(n5212), .A3(n5198), .A4(n5352), .Z(n5423) );
  ND3D0 U5318 ( .A1(n5278), .A2(n4144), .A3(n5448), .ZN(n5352) );
  OR3D0 U5319 ( .A1(n5449), .A2(n5450), .A3(n5192), .Z(n5198) );
  OAI211D0 U5320 ( .A1(n5450), .A2(n5192), .B(n4119), .C(n5451), .ZN(n5212) );
  NR2D0 U5321 ( .A1(n5449), .A2(n5360), .ZN(n5451) );
  OAI211D0 U5322 ( .A1(n3506), .A2(n3318), .B(n3397), .C(n5452), .ZN(n5360) );
  AN2D0 U5323 ( .A1(n3410), .A2(n3411), .Z(n5452) );
  OA21D0 U5324 ( .A1(n3498), .A2(n3365), .B(n3493), .Z(n3397) );
  OA31D0 U5325 ( .A1(n5453), .A2(n5454), .A3(n3373), .B(n5455), .Z(n3493) );
  OAI31D0 U5326 ( .A1(fifo_7_snoop[0]), .A2(fifo_7_snoop[2]), .A3(
        fifo_7_snoop[1]), .B(n5456), .ZN(n3373) );
  CKND0 U5327 ( .I(fifo_7_snoop[3]), .ZN(n5456) );
  CKND2D0 U5328 ( .A1(n3371), .A2(n3372), .ZN(n5453) );
  CKND0 U5329 ( .I(n3377), .ZN(n3498) );
  OAI31D0 U5330 ( .A1(n5457), .A2(n5458), .A3(n5459), .B(n5460), .ZN(n3377) );
  CKND0 U5331 ( .I(n3389), .ZN(n3506) );
  CKND2D0 U5332 ( .A1(n5461), .A2(n5462), .ZN(n3389) );
  OAI21D0 U5333 ( .A1(n4146), .A2(n5295), .B(n5448), .ZN(n5449) );
  INR3D0 U5334 ( .A1(n5463), .B1(n5464), .B2(n5465), .ZN(n5448) );
  OAI211D0 U5335 ( .A1(n3375), .A2(n3365), .B(n3492), .C(n5466), .ZN(n5192) );
  OA211D0 U5336 ( .A1(n3318), .A2(n5467), .B(n3511), .C(n3510), .Z(n5466) );
  NR2D0 U5337 ( .A1(n3382), .A2(n3384), .ZN(n5467) );
  CKND0 U5338 ( .I(n5468), .ZN(n3384) );
  CKND0 U5339 ( .I(n5469), .ZN(n3382) );
  OA31D0 U5340 ( .A1(n3371), .A2(n4014), .A3(n5454), .B(n5470), .Z(n3492) );
  CKND0 U5341 ( .I(n3372), .ZN(n4014) );
  OAI31D0 U5342 ( .A1(fifo_6_snoop[0]), .A2(fifo_6_snoop[2]), .A3(
        fifo_6_snoop[1]), .B(n5471), .ZN(n3371) );
  CKND0 U5343 ( .I(fifo_6_snoop[3]), .ZN(n5471) );
  AOI21D0 U5344 ( .A1(n5472), .A2(n5458), .B(n5473), .ZN(n3375) );
  AN4D0 U5345 ( .A1(n5348), .A2(n5349), .A3(n5320), .A4(n4150), .Z(n5302) );
  IND3D0 U5346 ( .A1(n5465), .B1(n5463), .B2(n5464), .ZN(n5320) );
  NR2D0 U5347 ( .A1(n5337), .A2(n4456), .ZN(n5464) );
  CKND2D0 U5348 ( .A1(n5465), .A2(n5463), .ZN(n5349) );
  OA21D0 U5349 ( .A1(n5231), .A2(n5238), .B(n4150), .Z(n5463) );
  NR2D0 U5350 ( .A1(n5308), .A2(n4457), .ZN(n5465) );
  ND3D0 U5351 ( .A1(n4151), .A2(n4150), .A3(n5232), .ZN(n5348) );
  CKND0 U5352 ( .I(n5238), .ZN(n5232) );
  OAI221D0 U5353 ( .A1(n3497), .A2(n3365), .B1(n3504), .B2(n3318), .C(n5474), 
        .ZN(n5238) );
  NR2D0 U5354 ( .A1(n3491), .A2(n3509), .ZN(n5474) );
  OAI22D0 U5355 ( .A1(n5475), .A2(n5476), .B1(n4479), .B2(n5231), .ZN(n3509)
         );
  OAI22D0 U5356 ( .A1(n5477), .A2(n5478), .B1(n5479), .B2(n3361), .ZN(n3491)
         );
  CKND0 U5357 ( .I(n5480), .ZN(n5477) );
  OA22D0 U5358 ( .A1(n5481), .A2(n5482), .B1(n5483), .B2(n5484), .Z(n3504) );
  OA22D0 U5359 ( .A1(n5485), .A2(n5486), .B1(n5487), .B2(n5488), .Z(n3497) );
  CKND0 U5360 ( .I(n3926), .ZN(n4098) );
  CKND0 U5361 ( .I(n5295), .ZN(n5278) );
  OAI211D0 U5362 ( .A1(n5489), .A2(n3318), .B(n3398), .C(n3391), .ZN(n5295) );
  CKND0 U5363 ( .I(n3415), .ZN(n3391) );
  CKND2D0 U5364 ( .A1(n5490), .A2(n5491), .ZN(n3415) );
  OA221D0 U5365 ( .A1(n5454), .A2(n3372), .B1(n3394), .B2(n3365), .C(n5492), 
        .Z(n3398) );
  AN2D0 U5366 ( .A1(n5493), .A2(n5494), .Z(n3394) );
  OAI31D0 U5367 ( .A1(fifo_5_snoop[0]), .A2(fifo_5_snoop[2]), .A3(
        fifo_5_snoop[1]), .B(n5495), .ZN(n3372) );
  CKND0 U5368 ( .I(fifo_5_snoop[3]), .ZN(n5495) );
  ND3D0 U5369 ( .A1(n5496), .A2(n3370), .A3(n3369), .ZN(n5454) );
  NR2D0 U5370 ( .A1(n3385), .A2(n3383), .ZN(n5489) );
  CKND0 U5371 ( .I(n5497), .ZN(n3383) );
  CKND0 U5372 ( .I(n5498), .ZN(n3385) );
  CKND0 U5373 ( .I(n5308), .ZN(n5303) );
  IND4D0 U5374 ( .A1(n3401), .B1(n3413), .B2(n5499), .B3(n3409), .ZN(n5308) );
  NR2D0 U5375 ( .A1(n3405), .A2(n3406), .ZN(n5499) );
  OAI211D0 U5376 ( .A1(n5500), .A2(n3365), .B(n3360), .C(n3496), .ZN(n3401) );
  ND3D0 U5377 ( .A1(n5501), .A2(n3361), .A3(n3359), .ZN(n3360) );
  NR2D0 U5378 ( .A1(n3503), .A2(n3502), .ZN(n5500) );
  CKND0 U5379 ( .I(n5337), .ZN(n5325) );
  IND4D0 U5380 ( .A1(n5502), .B1(n3392), .B2(n3393), .B3(n5503), .ZN(n5337) );
  OAI222D0 U5381 ( .A1(n5504), .A2(n3318), .B1(n3395), .B2(n3365), .C1(n5505), 
        .C2(n3370), .ZN(n5502) );
  CKND2D0 U5382 ( .A1(n4016), .A2(n5496), .ZN(n3370) );
  AOI22D0 U5383 ( .A1(n5506), .A2(n5507), .B1(n5508), .B2(n5509), .ZN(n3395)
         );
  CKND0 U5384 ( .I(n5510), .ZN(n5507) );
  CKND2D0 U5385 ( .A1(n3500), .A2(n5442), .ZN(n3318) );
  CKND0 U5386 ( .I(n3365), .ZN(n5442) );
  CKND2D0 U5387 ( .A1(n3369), .A2(n5511), .ZN(n3365) );
  CKND0 U5388 ( .I(n5505), .ZN(n3369) );
  IND3D0 U5389 ( .A1(n5501), .B1(n3361), .B2(n3359), .ZN(n5505) );
  CKND0 U5390 ( .I(n5479), .ZN(n3359) );
  OAI21D0 U5391 ( .A1(n3374), .A2(n4283), .B(n5441), .ZN(n5479) );
  IND2D0 U5392 ( .A1(n3894), .B1(n5496), .ZN(n5441) );
  OAI31D0 U5393 ( .A1(fifo_0_snoop[0]), .A2(fifo_0_snoop[2]), .A3(
        fifo_0_snoop[1]), .B(n5512), .ZN(n4283) );
  CKND0 U5394 ( .I(fifo_0_snoop[3]), .ZN(n5512) );
  CKND2D0 U5395 ( .A1(n5496), .A2(n4019), .ZN(n3361) );
  OA31D0 U5396 ( .A1(fifo_2_snoop[0]), .A2(fifo_2_snoop[2]), .A3(
        fifo_2_snoop[1]), .B(n5513), .Z(n4019) );
  CKND0 U5397 ( .I(fifo_2_snoop[3]), .ZN(n5513) );
  CKND0 U5398 ( .I(n3374), .ZN(n5496) );
  NR2D0 U5399 ( .A1(n4011), .A2(n3374), .ZN(n5501) );
  CKND2D0 U5400 ( .A1(n3282), .A2(n5514), .ZN(n3374) );
  AN4D0 U5401 ( .A1(n3366), .A2(n3496), .A3(n5478), .A4(n5480), .Z(n3282) );
  IND3D0 U5402 ( .A1(n5515), .B1(n5478), .B2(n5480), .ZN(n3496) );
  AN4D0 U5403 ( .A1(n5503), .A2(n5492), .A3(n5470), .A4(n5455), .Z(n3366) );
  ND4D0 U5404 ( .A1(n4028), .A2(n5516), .A3(n5517), .A4(n5518), .ZN(n5455) );
  OA31D0 U5405 ( .A1(fifo_7_snoop[4]), .A2(fifo_7_snoop[6]), .A3(
        fifo_7_snoop[5]), .B(n5519), .Z(n4028) );
  CKND0 U5406 ( .I(fifo_7_snoop[7]), .ZN(n5519) );
  ND3D0 U5407 ( .A1(n5516), .A2(n5518), .A3(n4034), .ZN(n5470) );
  CKND0 U5408 ( .I(n5517), .ZN(n4034) );
  OAI31D0 U5409 ( .A1(fifo_6_snoop[4]), .A2(fifo_6_snoop[6]), .A3(
        fifo_6_snoop[5]), .B(n5520), .ZN(n5517) );
  CKND0 U5410 ( .I(fifo_6_snoop[7]), .ZN(n5520) );
  CKND2D0 U5411 ( .A1(n4029), .A2(n5516), .ZN(n5492) );
  AN3D0 U5412 ( .A1(n5514), .A2(n5521), .A3(n5511), .Z(n5516) );
  CKND0 U5413 ( .I(n5518), .ZN(n4029) );
  OAI31D0 U5414 ( .A1(fifo_5_snoop[4]), .A2(fifo_5_snoop[6]), .A3(
        fifo_5_snoop[5]), .B(n5522), .ZN(n5518) );
  CKND0 U5415 ( .I(fifo_5_snoop[7]), .ZN(n5522) );
  IND2D0 U5416 ( .A1(n5521), .B1(n5511), .ZN(n5503) );
  AN3D0 U5417 ( .A1(n5478), .A2(n5480), .A3(n5515), .Z(n5511) );
  CKND2D0 U5418 ( .A1(n4038), .A2(n5514), .ZN(n5515) );
  OA31D0 U5419 ( .A1(fifo_3_snoop[4]), .A2(fifo_3_snoop[6]), .A3(
        fifo_3_snoop[5]), .B(n5523), .Z(n4038) );
  CKND0 U5420 ( .I(fifo_3_snoop[7]), .ZN(n5523) );
  OAI21D0 U5421 ( .A1(n4035), .A2(n4352), .B(n5514), .ZN(n5480) );
  CKND0 U5422 ( .I(n4036), .ZN(n4352) );
  OAI31D0 U5423 ( .A1(fifo_1_snoop[4]), .A2(fifo_1_snoop[6]), .A3(
        fifo_1_snoop[5]), .B(n5524), .ZN(n4036) );
  CKND0 U5424 ( .I(fifo_1_snoop[7]), .ZN(n5524) );
  CKND0 U5425 ( .I(n3903), .ZN(n4035) );
  OAI31D0 U5426 ( .A1(fifo_0_snoop[4]), .A2(fifo_0_snoop[6]), .A3(
        fifo_0_snoop[5]), .B(n5525), .ZN(n3903) );
  CKND0 U5427 ( .I(fifo_0_snoop[7]), .ZN(n5525) );
  CKND2D0 U5428 ( .A1(n4037), .A2(n5514), .ZN(n5478) );
  OA31D0 U5429 ( .A1(fifo_2_snoop[4]), .A2(fifo_2_snoop[6]), .A3(
        fifo_2_snoop[5]), .B(n5526), .Z(n4037) );
  CKND0 U5430 ( .I(fifo_2_snoop[7]), .ZN(n5526) );
  CKND2D0 U5431 ( .A1(n4033), .A2(n5514), .ZN(n5521) );
  CKND0 U5432 ( .I(n5440), .ZN(n5514) );
  CKND2D0 U5433 ( .A1(n3283), .A2(n5527), .ZN(n5440) );
  CKND0 U5434 ( .I(n5528), .ZN(n3283) );
  IND4D0 U5435 ( .A1(n5458), .B1(n5494), .B2(n5457), .B3(n5529), .ZN(n5528) );
  NR4D0 U5436 ( .A1(n5509), .A2(n5487), .A3(n3503), .A4(n5530), .ZN(n5529) );
  NR3D0 U5437 ( .A1(n5530), .A2(n5487), .A3(n5531), .ZN(n3503) );
  CKND0 U5438 ( .I(n5532), .ZN(n5509) );
  OR2D0 U5439 ( .A1(n4043), .A2(n5445), .Z(n5457) );
  OAI31D0 U5440 ( .A1(fifo_7_snoop[10]), .A2(fifo_7_snoop[9]), .A3(
        fifo_7_snoop[8]), .B(n5533), .ZN(n4043) );
  CKND0 U5441 ( .I(fifo_7_snoop[11]), .ZN(n5533) );
  ND3D0 U5442 ( .A1(n5534), .A2(n5532), .A3(n5508), .ZN(n5494) );
  NR2D0 U5443 ( .A1(n4302), .A2(n5445), .ZN(n5458) );
  OAI31D0 U5444 ( .A1(fifo_6_snoop[10]), .A2(fifo_6_snoop[9]), .A3(
        fifo_6_snoop[8]), .B(n5535), .ZN(n4302) );
  CKND0 U5445 ( .I(fifo_6_snoop[11]), .ZN(n5535) );
  OA31D0 U5446 ( .A1(fifo_4_snoop[4]), .A2(fifo_4_snoop[6]), .A3(
        fifo_4_snoop[5]), .B(n5536), .Z(n4033) );
  CKND0 U5447 ( .I(fifo_4_snoop[7]), .ZN(n5536) );
  OAI31D0 U5448 ( .A1(fifo_3_snoop[0]), .A2(fifo_3_snoop[2]), .A3(
        fifo_3_snoop[1]), .B(n5537), .ZN(n4011) );
  CKND0 U5449 ( .I(fifo_3_snoop[3]), .ZN(n5537) );
  CKND0 U5450 ( .I(n3381), .ZN(n3500) );
  CKND2D0 U5451 ( .A1(n5472), .A2(n5538), .ZN(n3381) );
  CKND0 U5452 ( .I(n5459), .ZN(n5472) );
  IND3D0 U5453 ( .A1(n5534), .B1(n5508), .B2(n5532), .ZN(n5459) );
  CKND2D0 U5454 ( .A1(n4053), .A2(n5527), .ZN(n5532) );
  OA31D0 U5455 ( .A1(fifo_4_snoop[10]), .A2(fifo_4_snoop[9]), .A3(
        fifo_4_snoop[8]), .B(n5539), .Z(n4053) );
  CKND0 U5456 ( .I(fifo_4_snoop[11]), .ZN(n5539) );
  INR3D0 U5457 ( .A1(n5531), .B1(n5530), .B2(n5487), .ZN(n5508) );
  AOI21D0 U5458 ( .A1(n4050), .A2(n3910), .B(n5445), .ZN(n5487) );
  OAI31D0 U5459 ( .A1(fifo_0_snoop[10]), .A2(fifo_0_snoop[9]), .A3(
        fifo_0_snoop[8]), .B(n5540), .ZN(n3910) );
  CKND0 U5460 ( .I(fifo_0_snoop[11]), .ZN(n5540) );
  OAI31D0 U5461 ( .A1(fifo_1_snoop[10]), .A2(fifo_1_snoop[9]), .A3(
        fifo_1_snoop[8]), .B(n5541), .ZN(n4050) );
  CKND0 U5462 ( .I(fifo_1_snoop[11]), .ZN(n5541) );
  CKND0 U5463 ( .I(n5488), .ZN(n5530) );
  CKND2D0 U5464 ( .A1(n4052), .A2(n5527), .ZN(n5488) );
  OA31D0 U5465 ( .A1(fifo_2_snoop[10]), .A2(fifo_2_snoop[9]), .A3(
        fifo_2_snoop[8]), .B(n5542), .Z(n4052) );
  CKND0 U5466 ( .I(fifo_2_snoop[11]), .ZN(n5542) );
  CKND2D0 U5467 ( .A1(n4051), .A2(n5527), .ZN(n5531) );
  CKND0 U5468 ( .I(n5445), .ZN(n5527) );
  CKND0 U5469 ( .I(n3961), .ZN(n4051) );
  OAI31D0 U5470 ( .A1(fifo_3_snoop[10]), .A2(fifo_3_snoop[9]), .A3(
        fifo_3_snoop[8]), .B(n5543), .ZN(n3961) );
  CKND0 U5471 ( .I(fifo_3_snoop[11]), .ZN(n5543) );
  NR2D0 U5472 ( .A1(n4045), .A2(n5445), .ZN(n5534) );
  CKND2D0 U5473 ( .A1(n3284), .A2(n5544), .ZN(n5445) );
  AN4D0 U5474 ( .A1(n5493), .A2(n5460), .A3(n5510), .A4(n5545), .Z(n3284) );
  NR4D0 U5475 ( .A1(n5485), .A2(n3502), .A3(n5473), .A4(n5546), .ZN(n5545) );
  INR2D0 U5476 ( .A1(n5538), .B1(n5547), .ZN(n5473) );
  NR3D0 U5477 ( .A1(n5546), .A2(n5485), .A3(n5548), .ZN(n3502) );
  ND4D0 U5478 ( .A1(n4060), .A2(n5538), .A3(n5544), .A4(n5547), .ZN(n5460) );
  CKND2D0 U5479 ( .A1(n4062), .A2(n5544), .ZN(n5547) );
  OA31D0 U5480 ( .A1(fifo_6_snoop[12]), .A2(fifo_6_snoop[14]), .A3(
        fifo_6_snoop[13]), .B(n5549), .Z(n4062) );
  CKND0 U5481 ( .I(fifo_6_snoop[15]), .ZN(n5549) );
  AN3D0 U5482 ( .A1(n5550), .A2(n5510), .A3(n5506), .Z(n5538) );
  OA31D0 U5483 ( .A1(fifo_7_snoop[12]), .A2(fifo_7_snoop[14]), .A3(
        fifo_7_snoop[13]), .B(n5551), .Z(n4060) );
  CKND0 U5484 ( .I(fifo_7_snoop[15]), .ZN(n5551) );
  IND3D0 U5485 ( .A1(n5550), .B1(n5506), .B2(n5510), .ZN(n5493) );
  CKND2D0 U5486 ( .A1(n4066), .A2(n5544), .ZN(n5510) );
  OA31D0 U5487 ( .A1(fifo_4_snoop[12]), .A2(fifo_4_snoop[14]), .A3(
        fifo_4_snoop[13]), .B(n5552), .Z(n4066) );
  CKND0 U5488 ( .I(fifo_4_snoop[15]), .ZN(n5552) );
  INR3D0 U5489 ( .A1(n5548), .B1(n5546), .B2(n5485), .ZN(n5506) );
  AOI21D0 U5490 ( .A1(n3916), .A2(n4068), .B(n5444), .ZN(n5485) );
  CKND0 U5491 ( .I(n5544), .ZN(n5444) );
  OAI31D0 U5492 ( .A1(fifo_1_snoop[12]), .A2(fifo_1_snoop[14]), .A3(
        fifo_1_snoop[13]), .B(n5553), .ZN(n4068) );
  CKND0 U5493 ( .I(fifo_1_snoop[15]), .ZN(n5553) );
  OAI31D0 U5494 ( .A1(fifo_0_snoop[12]), .A2(fifo_0_snoop[14]), .A3(
        fifo_0_snoop[13]), .B(n5554), .ZN(n3916) );
  CKND0 U5495 ( .I(fifo_0_snoop[15]), .ZN(n5554) );
  CKND0 U5496 ( .I(n5486), .ZN(n5546) );
  CKND2D0 U5497 ( .A1(n4069), .A2(n5544), .ZN(n5486) );
  OA31D0 U5498 ( .A1(fifo_2_snoop[12]), .A2(fifo_2_snoop[14]), .A3(
        fifo_2_snoop[13]), .B(n5555), .Z(n4069) );
  CKND0 U5499 ( .I(fifo_2_snoop[15]), .ZN(n5555) );
  CKND2D0 U5500 ( .A1(n4070), .A2(n5544), .ZN(n5548) );
  OA31D0 U5501 ( .A1(fifo_3_snoop[12]), .A2(fifo_3_snoop[14]), .A3(
        fifo_3_snoop[13]), .B(n5556), .Z(n4070) );
  CKND0 U5502 ( .I(fifo_3_snoop[15]), .ZN(n5556) );
  CKND2D0 U5503 ( .A1(n4065), .A2(n5544), .ZN(n5550) );
  NR2D0 U5504 ( .A1(n3320), .A2(n5447), .ZN(n5544) );
  ND4D0 U5505 ( .A1(n5498), .A2(n5468), .A3(n5557), .A4(n5558), .ZN(n3320) );
  INR4D0 U5506 ( .A1(n5461), .B1(n5483), .B2(n3406), .B3(n5559), .ZN(n5558) );
  INR3D0 U5507 ( .A1(n5560), .B1(n5559), .B2(n5483), .ZN(n3406) );
  ND4D0 U5508 ( .A1(n4326), .A2(n5561), .A3(n4073), .A4(n4074), .ZN(n5461) );
  CKND0 U5509 ( .I(n4077), .ZN(n4326) );
  OAI31D0 U5510 ( .A1(fifo_7_snoop[16]), .A2(fifo_7_snoop[18]), .A3(
        fifo_7_snoop[17]), .B(n5562), .ZN(n4077) );
  CKND0 U5511 ( .I(fifo_7_snoop[19]), .ZN(n5562) );
  ND3D0 U5512 ( .A1(n5561), .A2(n4074), .A3(n4076), .ZN(n5468) );
  CKND0 U5513 ( .I(n4073), .ZN(n4076) );
  OAI31D0 U5514 ( .A1(fifo_6_snoop[16]), .A2(fifo_6_snoop[18]), .A3(
        fifo_6_snoop[17]), .B(n5563), .ZN(n4073) );
  CKND0 U5515 ( .I(fifo_6_snoop[19]), .ZN(n5563) );
  CKND2D0 U5516 ( .A1(n5157), .A2(n5561), .ZN(n5498) );
  INR3D0 U5517 ( .A1(n5557), .B1(n3512), .B2(n5447), .ZN(n5561) );
  CKND0 U5518 ( .I(n4074), .ZN(n5157) );
  OAI31D0 U5519 ( .A1(fifo_5_snoop[16]), .A2(fifo_5_snoop[18]), .A3(
        fifo_5_snoop[17]), .B(n5564), .ZN(n4074) );
  CKND0 U5520 ( .I(fifo_5_snoop[19]), .ZN(n5564) );
  OA31D0 U5521 ( .A1(fifo_5_snoop[12]), .A2(fifo_5_snoop[14]), .A3(
        fifo_5_snoop[13]), .B(n5565), .Z(n4065) );
  CKND0 U5522 ( .I(fifo_5_snoop[15]), .ZN(n5565) );
  OAI31D0 U5523 ( .A1(fifo_5_snoop[10]), .A2(fifo_5_snoop[9]), .A3(
        fifo_5_snoop[8]), .B(n5566), .ZN(n4045) );
  CKND0 U5524 ( .I(fifo_5_snoop[11]), .ZN(n5566) );
  CKND0 U5525 ( .I(n3388), .ZN(n5504) );
  OAI22D0 U5526 ( .A1(n3513), .A2(n5567), .B1(n3512), .B2(n5557), .ZN(n3388)
         );
  CKND2D0 U5527 ( .A1(n4083), .A2(n5568), .ZN(n5557) );
  OA31D0 U5528 ( .A1(fifo_4_snoop[16]), .A2(fifo_4_snoop[18]), .A3(
        fifo_4_snoop[17]), .B(n5569), .Z(n4083) );
  CKND0 U5529 ( .I(fifo_4_snoop[19]), .ZN(n5569) );
  OR3D0 U5530 ( .A1(n5559), .A2(n5483), .A3(n5560), .Z(n3512) );
  NR2D0 U5531 ( .A1(n4004), .A2(n5447), .ZN(n5560) );
  OAI31D0 U5532 ( .A1(fifo_3_snoop[16]), .A2(fifo_3_snoop[18]), .A3(
        fifo_3_snoop[17]), .B(n5570), .ZN(n4004) );
  CKND0 U5533 ( .I(fifo_3_snoop[19]), .ZN(n5570) );
  AOI21D0 U5534 ( .A1(n3922), .A2(n4080), .B(n5447), .ZN(n5483) );
  CKND0 U5535 ( .I(n5568), .ZN(n5447) );
  OAI31D0 U5536 ( .A1(fifo_1_snoop[16]), .A2(fifo_1_snoop[18]), .A3(
        fifo_1_snoop[17]), .B(n5571), .ZN(n4080) );
  CKND0 U5537 ( .I(fifo_1_snoop[19]), .ZN(n5571) );
  OAI31D0 U5538 ( .A1(fifo_0_snoop[16]), .A2(fifo_0_snoop[18]), .A3(
        fifo_0_snoop[17]), .B(n5572), .ZN(n3922) );
  CKND0 U5539 ( .I(fifo_0_snoop[19]), .ZN(n5572) );
  CKND0 U5540 ( .I(n5484), .ZN(n5559) );
  CKND2D0 U5541 ( .A1(n4082), .A2(n5568), .ZN(n5484) );
  NR2D0 U5542 ( .A1(n3319), .A2(n5446), .ZN(n5568) );
  ND4D0 U5543 ( .A1(n5497), .A2(n5469), .A3(n5567), .A4(n5573), .ZN(n3319) );
  INR4D0 U5544 ( .A1(n5462), .B1(n5481), .B2(n3405), .B3(n5574), .ZN(n5573) );
  NR3D0 U5545 ( .A1(n5574), .A2(n5481), .A3(n5575), .ZN(n3405) );
  CKND0 U5546 ( .I(n5482), .ZN(n5574) );
  ND4D0 U5547 ( .A1(n4310), .A2(n5576), .A3(n5577), .A4(n5578), .ZN(n5462) );
  CKND0 U5548 ( .I(n4092), .ZN(n4310) );
  OAI31D0 U5549 ( .A1(fifo_7_snoop[20]), .A2(fifo_7_snoop[22]), .A3(
        fifo_7_snoop[21]), .B(n5579), .ZN(n4092) );
  CKND0 U5550 ( .I(fifo_7_snoop[23]), .ZN(n5579) );
  ND3D0 U5551 ( .A1(n5576), .A2(n5577), .A3(n4097), .ZN(n5469) );
  CKND0 U5552 ( .I(n5578), .ZN(n4097) );
  OAI31D0 U5553 ( .A1(fifo_6_snoop[20]), .A2(fifo_6_snoop[22]), .A3(
        fifo_6_snoop[21]), .B(n5580), .ZN(n5578) );
  CKND0 U5554 ( .I(fifo_6_snoop[23]), .ZN(n5580) );
  CKND2D0 U5555 ( .A1(n4087), .A2(n5576), .ZN(n5497) );
  INR3D0 U5556 ( .A1(n5567), .B1(n3513), .B2(n5446), .ZN(n5576) );
  CKND0 U5557 ( .I(n5577), .ZN(n4087) );
  OAI31D0 U5558 ( .A1(fifo_5_snoop[20]), .A2(fifo_5_snoop[22]), .A3(
        fifo_5_snoop[21]), .B(n5581), .ZN(n5577) );
  CKND0 U5559 ( .I(fifo_5_snoop[23]), .ZN(n5581) );
  OA31D0 U5560 ( .A1(fifo_2_snoop[16]), .A2(fifo_2_snoop[18]), .A3(
        fifo_2_snoop[17]), .B(n5582), .Z(n4082) );
  CKND0 U5561 ( .I(fifo_2_snoop[19]), .ZN(n5582) );
  CKND2D0 U5562 ( .A1(n4096), .A2(n5583), .ZN(n5567) );
  OA31D0 U5563 ( .A1(fifo_4_snoop[20]), .A2(fifo_4_snoop[22]), .A3(
        fifo_4_snoop[21]), .B(n5584), .Z(n4096) );
  CKND0 U5564 ( .I(fifo_4_snoop[23]), .ZN(n5584) );
  IND3D0 U5565 ( .A1(n5481), .B1(n5575), .B2(n5482), .ZN(n3513) );
  CKND2D0 U5566 ( .A1(n4100), .A2(n5583), .ZN(n5482) );
  OA31D0 U5567 ( .A1(fifo_2_snoop[20]), .A2(fifo_2_snoop[22]), .A3(
        fifo_2_snoop[21]), .B(n5585), .Z(n4100) );
  CKND0 U5568 ( .I(fifo_2_snoop[23]), .ZN(n5585) );
  CKND2D0 U5569 ( .A1(n4101), .A2(n5583), .ZN(n5575) );
  CKND0 U5570 ( .I(n5446), .ZN(n5583) );
  OA31D0 U5571 ( .A1(fifo_3_snoop[20]), .A2(fifo_3_snoop[22]), .A3(
        fifo_3_snoop[21]), .B(n5586), .Z(n4101) );
  CKND0 U5572 ( .I(fifo_3_snoop[23]), .ZN(n5586) );
  AOI21D0 U5573 ( .A1(n3926), .A2(n4099), .B(n5446), .ZN(n5481) );
  CKND2D0 U5574 ( .A1(n3358), .A2(n5587), .ZN(n5446) );
  AN4D0 U5575 ( .A1(n5490), .A2(n3413), .A3(n3392), .A4(n5588), .Z(n3358) );
  AN4D0 U5576 ( .A1(n5589), .A2(n5476), .A3(n3411), .A4(n3510), .Z(n5588) );
  ND3D0 U5577 ( .A1(n5590), .A2(n4114), .A3(n4106), .ZN(n3510) );
  CKND0 U5578 ( .I(n5591), .ZN(n4106) );
  ND4D0 U5579 ( .A1(n5427), .A2(n5590), .A3(n5591), .A4(n4114), .ZN(n3411) );
  OAI31D0 U5580 ( .A1(fifo_6_snoop[24]), .A2(fifo_6_snoop[26]), .A3(
        fifo_6_snoop[25]), .B(n5592), .ZN(n5591) );
  CKND0 U5581 ( .I(fifo_6_snoop[27]), .ZN(n5592) );
  CKND0 U5582 ( .I(n4107), .ZN(n5427) );
  OAI31D0 U5583 ( .A1(fifo_7_snoop[24]), .A2(fifo_7_snoop[26]), .A3(
        fifo_7_snoop[25]), .B(n5593), .ZN(n4107) );
  CKND0 U5584 ( .I(fifo_7_snoop[27]), .ZN(n5593) );
  ND3D0 U5585 ( .A1(n4115), .A2(n5587), .A3(n5594), .ZN(n3392) );
  ND3D0 U5586 ( .A1(n5476), .A2(n5589), .A3(n5595), .ZN(n3413) );
  CKND2D0 U5587 ( .A1(n5424), .A2(n5590), .ZN(n5490) );
  INR3D0 U5588 ( .A1(n5594), .B1(n5439), .B2(n4115), .ZN(n5590) );
  CKND0 U5589 ( .I(n4397), .ZN(n4115) );
  OAI31D0 U5590 ( .A1(fifo_4_snoop[24]), .A2(fifo_4_snoop[26]), .A3(
        fifo_4_snoop[25]), .B(n5596), .ZN(n4397) );
  CKND0 U5591 ( .I(fifo_4_snoop[27]), .ZN(n5596) );
  INR3D0 U5592 ( .A1(n5476), .B1(n5475), .B2(n5595), .ZN(n5594) );
  NR2D0 U5593 ( .A1(n4110), .A2(n5439), .ZN(n5595) );
  OAI31D0 U5594 ( .A1(fifo_3_snoop[24]), .A2(fifo_3_snoop[26]), .A3(
        fifo_3_snoop[25]), .B(n5597), .ZN(n4110) );
  CKND0 U5595 ( .I(fifo_3_snoop[27]), .ZN(n5597) );
  CKND0 U5596 ( .I(n5589), .ZN(n5475) );
  OAI21D0 U5597 ( .A1(n4112), .A2(n4111), .B(n5587), .ZN(n5589) );
  CKND0 U5598 ( .I(n5438), .ZN(n4111) );
  OAI31D0 U5599 ( .A1(fifo_1_snoop[24]), .A2(fifo_1_snoop[26]), .A3(
        fifo_1_snoop[25]), .B(n5598), .ZN(n5438) );
  CKND0 U5600 ( .I(fifo_1_snoop[27]), .ZN(n5598) );
  OA31D0 U5601 ( .A1(fifo_0_snoop[24]), .A2(fifo_0_snoop[26]), .A3(
        fifo_0_snoop[25]), .B(n5599), .Z(n4112) );
  CKND0 U5602 ( .I(fifo_0_snoop[27]), .ZN(n5599) );
  CKND2D0 U5603 ( .A1(n4113), .A2(n5587), .ZN(n5476) );
  CKND0 U5604 ( .I(n5439), .ZN(n5587) );
  ND4D0 U5605 ( .A1(n3511), .A2(n3410), .A3(n3409), .A4(n5600), .ZN(n5439) );
  AN3D0 U5606 ( .A1(n5491), .A2(n5601), .A3(n3393), .Z(n5600) );
  ND3D0 U5607 ( .A1(n5601), .A2(n4457), .A3(n4147), .ZN(n3393) );
  CKND2D0 U5608 ( .A1(n4144), .A2(n5602), .ZN(n5491) );
  CKND0 U5609 ( .I(n4146), .ZN(n4144) );
  CKND2D0 U5610 ( .A1(n4148), .A2(n5601), .ZN(n3409) );
  ND4D0 U5611 ( .A1(n4119), .A2(n5602), .A3(n5450), .A4(n4146), .ZN(n3410) );
  OA31D0 U5612 ( .A1(fifo_7_snoop[28]), .A2(fifo_7_snoop[30]), .A3(
        fifo_7_snoop[29]), .B(n5603), .Z(n4119) );
  CKND0 U5613 ( .I(fifo_7_snoop[31]), .ZN(n5603) );
  ND3D0 U5614 ( .A1(n5602), .A2(n4146), .A3(n4121), .ZN(n3511) );
  CKND0 U5615 ( .I(n5450), .ZN(n4121) );
  OAI31D0 U5616 ( .A1(fifo_6_snoop[28]), .A2(fifo_6_snoop[30]), .A3(
        fifo_6_snoop[29]), .B(n5604), .ZN(n5450) );
  CKND0 U5617 ( .I(fifo_6_snoop[31]), .ZN(n5604) );
  OAI31D0 U5618 ( .A1(fifo_5_snoop[28]), .A2(fifo_5_snoop[30]), .A3(
        fifo_5_snoop[29]), .B(n5605), .ZN(n4146) );
  CKND0 U5619 ( .I(fifo_5_snoop[31]), .ZN(n5605) );
  INR3D0 U5620 ( .A1(n5601), .B1(n4148), .B2(n4147), .ZN(n5602) );
  CKND0 U5621 ( .I(n4456), .ZN(n4147) );
  OAI31D0 U5622 ( .A1(fifo_4_snoop[28]), .A2(fifo_4_snoop[30]), .A3(
        fifo_4_snoop[29]), .B(n5606), .ZN(n4456) );
  CKND0 U5623 ( .I(fifo_4_snoop[31]), .ZN(n5606) );
  CKND0 U5624 ( .I(n4457), .ZN(n4148) );
  OAI31D0 U5625 ( .A1(fifo_3_snoop[28]), .A2(fifo_3_snoop[30]), .A3(
        fifo_3_snoop[29]), .B(n5607), .ZN(n4457) );
  CKND0 U5626 ( .I(fifo_3_snoop[31]), .ZN(n5607) );
  NR2D0 U5627 ( .A1(n4479), .A2(n4151), .ZN(n5601) );
  CKND0 U5628 ( .I(n5231), .ZN(n4151) );
  OAI31D0 U5629 ( .A1(fifo_2_snoop[28]), .A2(fifo_2_snoop[30]), .A3(
        fifo_2_snoop[29]), .B(n5608), .ZN(n5231) );
  CKND0 U5630 ( .I(fifo_2_snoop[31]), .ZN(n5608) );
  CKND2D0 U5631 ( .A1(n4150), .A2(n4149), .ZN(n4479) );
  OAI31D0 U5632 ( .A1(fifo_1_snoop[28]), .A2(fifo_1_snoop[30]), .A3(
        fifo_1_snoop[29]), .B(n5609), .ZN(n4149) );
  CKND0 U5633 ( .I(fifo_1_snoop[31]), .ZN(n5609) );
  OAI31D0 U5634 ( .A1(fifo_0_snoop[28]), .A2(fifo_0_snoop[30]), .A3(
        fifo_0_snoop[29]), .B(n5610), .ZN(n4150) );
  CKND0 U5635 ( .I(fifo_0_snoop[31]), .ZN(n5610) );
  OA31D0 U5636 ( .A1(fifo_2_snoop[24]), .A2(fifo_2_snoop[26]), .A3(
        fifo_2_snoop[25]), .B(n5611), .Z(n4113) );
  CKND0 U5637 ( .I(fifo_2_snoop[27]), .ZN(n5611) );
  CKND0 U5638 ( .I(n4114), .ZN(n5424) );
  OAI31D0 U5639 ( .A1(fifo_5_snoop[24]), .A2(fifo_5_snoop[26]), .A3(
        fifo_5_snoop[25]), .B(n5612), .ZN(n4114) );
  CKND0 U5640 ( .I(fifo_5_snoop[27]), .ZN(n5612) );
  OAI31D0 U5641 ( .A1(fifo_1_snoop[20]), .A2(fifo_1_snoop[22]), .A3(
        fifo_1_snoop[21]), .B(n5613), .ZN(n4099) );
  CKND0 U5642 ( .I(fifo_1_snoop[23]), .ZN(n5613) );
  OAI31D0 U5643 ( .A1(fifo_0_snoop[20]), .A2(fifo_0_snoop[22]), .A3(
        fifo_0_snoop[21]), .B(n5614), .ZN(n3926) );
  CKND0 U5644 ( .I(fifo_0_snoop[23]), .ZN(n5614) );
  OA31D0 U5645 ( .A1(fifo_4_snoop[0]), .A2(fifo_4_snoop[2]), .A3(
        fifo_4_snoop[1]), .B(n5615), .Z(n4016) );
  CKND0 U5646 ( .I(fifo_4_snoop[3]), .ZN(n5615) );
  OAI31D0 U5647 ( .A1(fifo_1_snoop[0]), .A2(fifo_1_snoop[2]), .A3(
        fifo_1_snoop[1]), .B(n5616), .ZN(n3894) );
  CKND0 U5648 ( .I(fifo_1_snoop[3]), .ZN(n5616) );
endmodule

