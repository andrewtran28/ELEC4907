
module crossbar_0 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_1 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_2 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_3 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_4 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_5 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_6 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_7 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_8 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_9 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_10 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_11 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_12 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_13 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_14 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_15 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_16 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_17 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_18 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module crossbar_19 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  MUX2ND0 U1 ( .I0(n1), .I1(n2), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n3), .I1(n4), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n5), .I1(n6), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n7), .I1(n8), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n9), .I1(n10), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n13), .I1(n14), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n15), .I1(n16), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n17), .I1(n18), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n19), .I1(n20), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n21), .I1(n22), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n23), .I1(n24), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n25), .I1(n26), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n27), .I1(n28), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n29), .I1(n30), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n31), .I1(n32), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n33), .I1(n34), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n35), .I1(n36), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n37), .I1(n38), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n39), .I1(n40), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n2), .I1(n1), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n1) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n2) );
  MUX2ND0 U24 ( .I0(n4), .I1(n3), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n3) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n4) );
  MUX2ND0 U27 ( .I0(n6), .I1(n5), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n5) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n6) );
  MUX2ND0 U30 ( .I0(n8), .I1(n7), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n7) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n8) );
  MUX2ND0 U33 ( .I0(n10), .I1(n9), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n9) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n10) );
  MUX2ND0 U36 ( .I0(n12), .I1(n11), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n11) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n12) );
  MUX2ND0 U39 ( .I0(n14), .I1(n13), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n13) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n14) );
  MUX2ND0 U42 ( .I0(n16), .I1(n15), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n15) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n16) );
  MUX2ND0 U45 ( .I0(n18), .I1(n17), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n17) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n18) );
  MUX2ND0 U48 ( .I0(n20), .I1(n19), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n19) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n20) );
  MUX2ND0 U51 ( .I0(n22), .I1(n21), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n21) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n22) );
  MUX2ND0 U54 ( .I0(n24), .I1(n23), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n23) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n24) );
  MUX2ND0 U57 ( .I0(n26), .I1(n25), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n25) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n26) );
  MUX2ND0 U60 ( .I0(n28), .I1(n27), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n27) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n28) );
  MUX2ND0 U63 ( .I0(n30), .I1(n29), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n29) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n30) );
  MUX2ND0 U66 ( .I0(n32), .I1(n31), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n31) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n32) );
  MUX2ND0 U69 ( .I0(n34), .I1(n33), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n33) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n34) );
  MUX2ND0 U72 ( .I0(n36), .I1(n35), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n35) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n36) );
  MUX2ND0 U75 ( .I0(n38), .I1(n37), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n37) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n38) );
  MUX2ND0 U78 ( .I0(n40), .I1(n39), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n39) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n40) );
endmodule


module benes ( in_input, in_control, port_en_n, out_output, clk, rst );
  input [127:0] in_input;
  input [19:0] in_control;
  input [7:0] port_en_n;
  output [159:0] out_output;
  input clk, rst;
  wire   \*Logic1* , \in_upper_00[3] , \in_lower_00[3] , \in_upper_01[3] ,
         \in_lower_01[3] , in_upper_02_3, \in_lower_02[3] , \in_upper_03[3] ,
         \stage_0_output[7][19] , \stage_0_output[7][18] ,
         \stage_0_output[7][17] , \stage_0_output[7][16] ,
         \stage_0_output[7][15] , \stage_0_output[7][14] ,
         \stage_0_output[7][13] , \stage_0_output[7][12] ,
         \stage_0_output[7][11] , \stage_0_output[7][10] ,
         \stage_0_output[7][9] , \stage_0_output[7][8] ,
         \stage_0_output[7][7] , \stage_0_output[7][6] ,
         \stage_0_output[7][5] , \stage_0_output[7][4] ,
         \stage_0_output[7][3] , \stage_0_output[7][2] ,
         \stage_0_output[7][1] , \stage_0_output[7][0] ,
         \stage_0_output[6][19] , \stage_0_output[6][18] ,
         \stage_0_output[6][17] , \stage_0_output[6][16] ,
         \stage_0_output[6][15] , \stage_0_output[6][14] ,
         \stage_0_output[6][13] , \stage_0_output[6][12] ,
         \stage_0_output[6][11] , \stage_0_output[6][10] ,
         \stage_0_output[6][9] , \stage_0_output[6][8] ,
         \stage_0_output[6][7] , \stage_0_output[6][6] ,
         \stage_0_output[6][5] , \stage_0_output[6][4] ,
         \stage_0_output[6][3] , \stage_0_output[6][2] ,
         \stage_0_output[6][1] , \stage_0_output[6][0] ,
         \stage_0_output[5][19] , \stage_0_output[5][18] ,
         \stage_0_output[5][17] , \stage_0_output[5][16] ,
         \stage_0_output[5][15] , \stage_0_output[5][14] ,
         \stage_0_output[5][13] , \stage_0_output[5][12] ,
         \stage_0_output[5][11] , \stage_0_output[5][10] ,
         \stage_0_output[5][9] , \stage_0_output[5][8] ,
         \stage_0_output[5][7] , \stage_0_output[5][6] ,
         \stage_0_output[5][5] , \stage_0_output[5][4] ,
         \stage_0_output[5][3] , \stage_0_output[5][2] ,
         \stage_0_output[5][1] , \stage_0_output[5][0] ,
         \stage_0_output[4][19] , \stage_0_output[4][18] ,
         \stage_0_output[4][17] , \stage_0_output[4][16] ,
         \stage_0_output[4][15] , \stage_0_output[4][14] ,
         \stage_0_output[4][13] , \stage_0_output[4][12] ,
         \stage_0_output[4][11] , \stage_0_output[4][10] ,
         \stage_0_output[4][9] , \stage_0_output[4][8] ,
         \stage_0_output[4][7] , \stage_0_output[4][6] ,
         \stage_0_output[4][5] , \stage_0_output[4][4] ,
         \stage_0_output[4][3] , \stage_0_output[4][2] ,
         \stage_0_output[4][1] , \stage_0_output[4][0] ,
         \stage_0_output[3][19] , \stage_0_output[3][18] ,
         \stage_0_output[3][17] , \stage_0_output[3][16] ,
         \stage_0_output[3][15] , \stage_0_output[3][14] ,
         \stage_0_output[3][13] , \stage_0_output[3][12] ,
         \stage_0_output[3][11] , \stage_0_output[3][10] ,
         \stage_0_output[3][9] , \stage_0_output[3][8] ,
         \stage_0_output[3][7] , \stage_0_output[3][6] ,
         \stage_0_output[3][5] , \stage_0_output[3][4] ,
         \stage_0_output[3][3] , \stage_0_output[3][2] ,
         \stage_0_output[3][1] , \stage_0_output[3][0] ,
         \stage_0_output[2][19] , \stage_0_output[2][18] ,
         \stage_0_output[2][17] , \stage_0_output[2][16] ,
         \stage_0_output[2][15] , \stage_0_output[2][14] ,
         \stage_0_output[2][13] , \stage_0_output[2][12] ,
         \stage_0_output[2][11] , \stage_0_output[2][10] ,
         \stage_0_output[2][9] , \stage_0_output[2][8] ,
         \stage_0_output[2][7] , \stage_0_output[2][6] ,
         \stage_0_output[2][5] , \stage_0_output[2][4] ,
         \stage_0_output[2][3] , \stage_0_output[2][2] ,
         \stage_0_output[2][1] , \stage_0_output[2][0] ,
         \stage_0_output[1][19] , \stage_0_output[1][18] ,
         \stage_0_output[1][17] , \stage_0_output[1][16] ,
         \stage_0_output[1][15] , \stage_0_output[1][14] ,
         \stage_0_output[1][13] , \stage_0_output[1][12] ,
         \stage_0_output[1][11] , \stage_0_output[1][10] ,
         \stage_0_output[1][9] , \stage_0_output[1][8] ,
         \stage_0_output[1][7] , \stage_0_output[1][6] ,
         \stage_0_output[1][5] , \stage_0_output[1][4] ,
         \stage_0_output[1][3] , \stage_0_output[1][2] ,
         \stage_0_output[1][1] , \stage_0_output[1][0] ,
         \stage_0_output[0][19] , \stage_0_output[0][18] ,
         \stage_0_output[0][17] , \stage_0_output[0][16] ,
         \stage_0_output[0][15] , \stage_0_output[0][14] ,
         \stage_0_output[0][13] , \stage_0_output[0][12] ,
         \stage_0_output[0][11] , \stage_0_output[0][10] ,
         \stage_0_output[0][9] , \stage_0_output[0][8] ,
         \stage_0_output[0][7] , \stage_0_output[0][6] ,
         \stage_0_output[0][5] , \stage_0_output[0][4] ,
         \stage_0_output[0][3] , \stage_0_output[0][2] ,
         \stage_0_output[0][1] , \stage_0_output[0][0] ,
         \stage_0_retimer[7][19] , \stage_0_retimer[7][18] ,
         \stage_0_retimer[7][17] , \stage_0_retimer[7][16] ,
         \stage_0_retimer[7][15] , \stage_0_retimer[7][14] ,
         \stage_0_retimer[7][13] , \stage_0_retimer[7][12] ,
         \stage_0_retimer[7][11] , \stage_0_retimer[7][10] ,
         \stage_0_retimer[7][9] , \stage_0_retimer[7][8] ,
         \stage_0_retimer[7][7] , \stage_0_retimer[7][6] ,
         \stage_0_retimer[7][5] , \stage_0_retimer[7][4] ,
         \stage_0_retimer[7][3] , \stage_0_retimer[7][2] ,
         \stage_0_retimer[7][1] , \stage_0_retimer[7][0] ,
         \stage_0_retimer[6][19] , \stage_0_retimer[6][18] ,
         \stage_0_retimer[6][17] , \stage_0_retimer[6][16] ,
         \stage_0_retimer[6][15] , \stage_0_retimer[6][14] ,
         \stage_0_retimer[6][13] , \stage_0_retimer[6][12] ,
         \stage_0_retimer[6][11] , \stage_0_retimer[6][10] ,
         \stage_0_retimer[6][9] , \stage_0_retimer[6][8] ,
         \stage_0_retimer[6][7] , \stage_0_retimer[6][6] ,
         \stage_0_retimer[6][5] , \stage_0_retimer[6][4] ,
         \stage_0_retimer[6][3] , \stage_0_retimer[6][2] ,
         \stage_0_retimer[6][1] , \stage_0_retimer[6][0] ,
         \stage_0_retimer[5][19] , \stage_0_retimer[5][18] ,
         \stage_0_retimer[5][17] , \stage_0_retimer[5][16] ,
         \stage_0_retimer[5][15] , \stage_0_retimer[5][14] ,
         \stage_0_retimer[5][13] , \stage_0_retimer[5][12] ,
         \stage_0_retimer[5][11] , \stage_0_retimer[5][10] ,
         \stage_0_retimer[5][9] , \stage_0_retimer[5][8] ,
         \stage_0_retimer[5][7] , \stage_0_retimer[5][6] ,
         \stage_0_retimer[5][5] , \stage_0_retimer[5][4] ,
         \stage_0_retimer[5][3] , \stage_0_retimer[5][2] ,
         \stage_0_retimer[5][1] , \stage_0_retimer[5][0] ,
         \stage_0_retimer[4][19] , \stage_0_retimer[4][18] ,
         \stage_0_retimer[4][17] , \stage_0_retimer[4][16] ,
         \stage_0_retimer[4][15] , \stage_0_retimer[4][14] ,
         \stage_0_retimer[4][13] , \stage_0_retimer[4][12] ,
         \stage_0_retimer[4][11] , \stage_0_retimer[4][10] ,
         \stage_0_retimer[4][9] , \stage_0_retimer[4][8] ,
         \stage_0_retimer[4][7] , \stage_0_retimer[4][6] ,
         \stage_0_retimer[4][5] , \stage_0_retimer[4][4] ,
         \stage_0_retimer[4][3] , \stage_0_retimer[4][2] ,
         \stage_0_retimer[4][1] , \stage_0_retimer[4][0] ,
         \stage_0_retimer[3][19] , \stage_0_retimer[3][18] ,
         \stage_0_retimer[3][17] , \stage_0_retimer[3][16] ,
         \stage_0_retimer[3][15] , \stage_0_retimer[3][14] ,
         \stage_0_retimer[3][13] , \stage_0_retimer[3][12] ,
         \stage_0_retimer[3][11] , \stage_0_retimer[3][10] ,
         \stage_0_retimer[3][9] , \stage_0_retimer[3][8] ,
         \stage_0_retimer[3][7] , \stage_0_retimer[3][6] ,
         \stage_0_retimer[3][5] , \stage_0_retimer[3][4] ,
         \stage_0_retimer[3][3] , \stage_0_retimer[3][2] ,
         \stage_0_retimer[3][1] , \stage_0_retimer[3][0] ,
         \stage_0_retimer[2][19] , \stage_0_retimer[2][18] ,
         \stage_0_retimer[2][17] , \stage_0_retimer[2][16] ,
         \stage_0_retimer[2][15] , \stage_0_retimer[2][14] ,
         \stage_0_retimer[2][13] , \stage_0_retimer[2][12] ,
         \stage_0_retimer[2][11] , \stage_0_retimer[2][10] ,
         \stage_0_retimer[2][9] , \stage_0_retimer[2][8] ,
         \stage_0_retimer[2][7] , \stage_0_retimer[2][6] ,
         \stage_0_retimer[2][5] , \stage_0_retimer[2][4] ,
         \stage_0_retimer[2][3] , \stage_0_retimer[2][2] ,
         \stage_0_retimer[2][1] , \stage_0_retimer[2][0] ,
         \stage_0_retimer[1][19] , \stage_0_retimer[1][18] ,
         \stage_0_retimer[1][17] , \stage_0_retimer[1][16] ,
         \stage_0_retimer[1][15] , \stage_0_retimer[1][14] ,
         \stage_0_retimer[1][13] , \stage_0_retimer[1][12] ,
         \stage_0_retimer[1][11] , \stage_0_retimer[1][10] ,
         \stage_0_retimer[1][9] , \stage_0_retimer[1][8] ,
         \stage_0_retimer[1][7] , \stage_0_retimer[1][6] ,
         \stage_0_retimer[1][5] , \stage_0_retimer[1][4] ,
         \stage_0_retimer[1][3] , \stage_0_retimer[1][2] ,
         \stage_0_retimer[1][1] , \stage_0_retimer[1][0] ,
         \stage_0_retimer[0][19] , \stage_0_retimer[0][18] ,
         \stage_0_retimer[0][17] , \stage_0_retimer[0][16] ,
         \stage_0_retimer[0][15] , \stage_0_retimer[0][14] ,
         \stage_0_retimer[0][13] , \stage_0_retimer[0][12] ,
         \stage_0_retimer[0][11] , \stage_0_retimer[0][10] ,
         \stage_0_retimer[0][9] , \stage_0_retimer[0][8] ,
         \stage_0_retimer[0][7] , \stage_0_retimer[0][6] ,
         \stage_0_retimer[0][5] , \stage_0_retimer[0][4] ,
         \stage_0_retimer[0][3] , \stage_0_retimer[0][2] ,
         \stage_0_retimer[0][1] , \stage_0_retimer[0][0] ,
         \stage_1_output[7][19] , \stage_1_output[7][18] ,
         \stage_1_output[7][17] , \stage_1_output[7][16] ,
         \stage_1_output[7][15] , \stage_1_output[7][14] ,
         \stage_1_output[7][13] , \stage_1_output[7][12] ,
         \stage_1_output[7][11] , \stage_1_output[7][10] ,
         \stage_1_output[7][9] , \stage_1_output[7][8] ,
         \stage_1_output[7][7] , \stage_1_output[7][6] ,
         \stage_1_output[7][5] , \stage_1_output[7][4] ,
         \stage_1_output[7][3] , \stage_1_output[7][2] ,
         \stage_1_output[7][1] , \stage_1_output[7][0] ,
         \stage_1_output[6][19] , \stage_1_output[6][18] ,
         \stage_1_output[6][17] , \stage_1_output[6][16] ,
         \stage_1_output[6][15] , \stage_1_output[6][14] ,
         \stage_1_output[6][13] , \stage_1_output[6][12] ,
         \stage_1_output[6][11] , \stage_1_output[6][10] ,
         \stage_1_output[6][9] , \stage_1_output[6][8] ,
         \stage_1_output[6][7] , \stage_1_output[6][6] ,
         \stage_1_output[6][5] , \stage_1_output[6][4] ,
         \stage_1_output[6][3] , \stage_1_output[6][2] ,
         \stage_1_output[6][1] , \stage_1_output[6][0] ,
         \stage_1_output[5][19] , \stage_1_output[5][18] ,
         \stage_1_output[5][17] , \stage_1_output[5][16] ,
         \stage_1_output[5][15] , \stage_1_output[5][14] ,
         \stage_1_output[5][13] , \stage_1_output[5][12] ,
         \stage_1_output[5][11] , \stage_1_output[5][10] ,
         \stage_1_output[5][9] , \stage_1_output[5][8] ,
         \stage_1_output[5][7] , \stage_1_output[5][6] ,
         \stage_1_output[5][5] , \stage_1_output[5][4] ,
         \stage_1_output[5][3] , \stage_1_output[5][2] ,
         \stage_1_output[5][1] , \stage_1_output[5][0] ,
         \stage_1_output[4][19] , \stage_1_output[4][18] ,
         \stage_1_output[4][17] , \stage_1_output[4][16] ,
         \stage_1_output[4][15] , \stage_1_output[4][14] ,
         \stage_1_output[4][13] , \stage_1_output[4][12] ,
         \stage_1_output[4][11] , \stage_1_output[4][10] ,
         \stage_1_output[4][9] , \stage_1_output[4][8] ,
         \stage_1_output[4][7] , \stage_1_output[4][6] ,
         \stage_1_output[4][5] , \stage_1_output[4][4] ,
         \stage_1_output[4][3] , \stage_1_output[4][2] ,
         \stage_1_output[4][1] , \stage_1_output[4][0] ,
         \stage_1_output[3][19] , \stage_1_output[3][18] ,
         \stage_1_output[3][17] , \stage_1_output[3][16] ,
         \stage_1_output[3][15] , \stage_1_output[3][14] ,
         \stage_1_output[3][13] , \stage_1_output[3][12] ,
         \stage_1_output[3][11] , \stage_1_output[3][10] ,
         \stage_1_output[3][9] , \stage_1_output[3][8] ,
         \stage_1_output[3][7] , \stage_1_output[3][6] ,
         \stage_1_output[3][5] , \stage_1_output[3][4] ,
         \stage_1_output[3][3] , \stage_1_output[3][2] ,
         \stage_1_output[3][1] , \stage_1_output[3][0] ,
         \stage_1_output[2][19] , \stage_1_output[2][18] ,
         \stage_1_output[2][17] , \stage_1_output[2][16] ,
         \stage_1_output[2][15] , \stage_1_output[2][14] ,
         \stage_1_output[2][13] , \stage_1_output[2][12] ,
         \stage_1_output[2][11] , \stage_1_output[2][10] ,
         \stage_1_output[2][9] , \stage_1_output[2][8] ,
         \stage_1_output[2][7] , \stage_1_output[2][6] ,
         \stage_1_output[2][5] , \stage_1_output[2][4] ,
         \stage_1_output[2][3] , \stage_1_output[2][2] ,
         \stage_1_output[2][1] , \stage_1_output[2][0] ,
         \stage_1_output[1][19] , \stage_1_output[1][18] ,
         \stage_1_output[1][17] , \stage_1_output[1][16] ,
         \stage_1_output[1][15] , \stage_1_output[1][14] ,
         \stage_1_output[1][13] , \stage_1_output[1][12] ,
         \stage_1_output[1][11] , \stage_1_output[1][10] ,
         \stage_1_output[1][9] , \stage_1_output[1][8] ,
         \stage_1_output[1][7] , \stage_1_output[1][6] ,
         \stage_1_output[1][5] , \stage_1_output[1][4] ,
         \stage_1_output[1][3] , \stage_1_output[1][2] ,
         \stage_1_output[1][1] , \stage_1_output[1][0] ,
         \stage_1_output[0][19] , \stage_1_output[0][18] ,
         \stage_1_output[0][17] , \stage_1_output[0][16] ,
         \stage_1_output[0][15] , \stage_1_output[0][14] ,
         \stage_1_output[0][13] , \stage_1_output[0][12] ,
         \stage_1_output[0][11] , \stage_1_output[0][10] ,
         \stage_1_output[0][9] , \stage_1_output[0][8] ,
         \stage_1_output[0][7] , \stage_1_output[0][6] ,
         \stage_1_output[0][5] , \stage_1_output[0][4] ,
         \stage_1_output[0][3] , \stage_1_output[0][2] ,
         \stage_1_output[0][1] , \stage_1_output[0][0] ,
         \stage_1_retimer[7][19] , \stage_1_retimer[7][18] ,
         \stage_1_retimer[7][17] , \stage_1_retimer[7][16] ,
         \stage_1_retimer[7][15] , \stage_1_retimer[7][14] ,
         \stage_1_retimer[7][13] , \stage_1_retimer[7][12] ,
         \stage_1_retimer[7][11] , \stage_1_retimer[7][10] ,
         \stage_1_retimer[7][9] , \stage_1_retimer[7][8] ,
         \stage_1_retimer[7][7] , \stage_1_retimer[7][6] ,
         \stage_1_retimer[7][5] , \stage_1_retimer[7][4] ,
         \stage_1_retimer[7][3] , \stage_1_retimer[7][2] ,
         \stage_1_retimer[7][1] , \stage_1_retimer[7][0] ,
         \stage_1_retimer[6][19] , \stage_1_retimer[6][18] ,
         \stage_1_retimer[6][17] , \stage_1_retimer[6][16] ,
         \stage_1_retimer[6][15] , \stage_1_retimer[6][14] ,
         \stage_1_retimer[6][13] , \stage_1_retimer[6][12] ,
         \stage_1_retimer[6][11] , \stage_1_retimer[6][10] ,
         \stage_1_retimer[6][9] , \stage_1_retimer[6][8] ,
         \stage_1_retimer[6][7] , \stage_1_retimer[6][6] ,
         \stage_1_retimer[6][5] , \stage_1_retimer[6][4] ,
         \stage_1_retimer[6][3] , \stage_1_retimer[6][2] ,
         \stage_1_retimer[6][1] , \stage_1_retimer[6][0] ,
         \stage_1_retimer[5][19] , \stage_1_retimer[5][18] ,
         \stage_1_retimer[5][17] , \stage_1_retimer[5][16] ,
         \stage_1_retimer[5][15] , \stage_1_retimer[5][14] ,
         \stage_1_retimer[5][13] , \stage_1_retimer[5][12] ,
         \stage_1_retimer[5][11] , \stage_1_retimer[5][10] ,
         \stage_1_retimer[5][9] , \stage_1_retimer[5][8] ,
         \stage_1_retimer[5][7] , \stage_1_retimer[5][6] ,
         \stage_1_retimer[5][5] , \stage_1_retimer[5][4] ,
         \stage_1_retimer[5][3] , \stage_1_retimer[5][2] ,
         \stage_1_retimer[5][1] , \stage_1_retimer[5][0] ,
         \stage_1_retimer[4][19] , \stage_1_retimer[4][18] ,
         \stage_1_retimer[4][17] , \stage_1_retimer[4][16] ,
         \stage_1_retimer[4][15] , \stage_1_retimer[4][14] ,
         \stage_1_retimer[4][13] , \stage_1_retimer[4][12] ,
         \stage_1_retimer[4][11] , \stage_1_retimer[4][10] ,
         \stage_1_retimer[4][9] , \stage_1_retimer[4][8] ,
         \stage_1_retimer[4][7] , \stage_1_retimer[4][6] ,
         \stage_1_retimer[4][5] , \stage_1_retimer[4][4] ,
         \stage_1_retimer[4][3] , \stage_1_retimer[4][2] ,
         \stage_1_retimer[4][1] , \stage_1_retimer[4][0] ,
         \stage_1_retimer[3][19] , \stage_1_retimer[3][18] ,
         \stage_1_retimer[3][17] , \stage_1_retimer[3][16] ,
         \stage_1_retimer[3][15] , \stage_1_retimer[3][14] ,
         \stage_1_retimer[3][13] , \stage_1_retimer[3][12] ,
         \stage_1_retimer[3][11] , \stage_1_retimer[3][10] ,
         \stage_1_retimer[3][9] , \stage_1_retimer[3][8] ,
         \stage_1_retimer[3][7] , \stage_1_retimer[3][6] ,
         \stage_1_retimer[3][5] , \stage_1_retimer[3][4] ,
         \stage_1_retimer[3][3] , \stage_1_retimer[3][2] ,
         \stage_1_retimer[3][1] , \stage_1_retimer[3][0] ,
         \stage_1_retimer[2][19] , \stage_1_retimer[2][18] ,
         \stage_1_retimer[2][17] , \stage_1_retimer[2][16] ,
         \stage_1_retimer[2][15] , \stage_1_retimer[2][14] ,
         \stage_1_retimer[2][13] , \stage_1_retimer[2][12] ,
         \stage_1_retimer[2][11] , \stage_1_retimer[2][10] ,
         \stage_1_retimer[2][9] , \stage_1_retimer[2][8] ,
         \stage_1_retimer[2][7] , \stage_1_retimer[2][6] ,
         \stage_1_retimer[2][5] , \stage_1_retimer[2][4] ,
         \stage_1_retimer[2][3] , \stage_1_retimer[2][2] ,
         \stage_1_retimer[2][1] , \stage_1_retimer[2][0] ,
         \stage_1_retimer[1][19] , \stage_1_retimer[1][18] ,
         \stage_1_retimer[1][17] , \stage_1_retimer[1][16] ,
         \stage_1_retimer[1][15] , \stage_1_retimer[1][14] ,
         \stage_1_retimer[1][13] , \stage_1_retimer[1][12] ,
         \stage_1_retimer[1][11] , \stage_1_retimer[1][10] ,
         \stage_1_retimer[1][9] , \stage_1_retimer[1][8] ,
         \stage_1_retimer[1][7] , \stage_1_retimer[1][6] ,
         \stage_1_retimer[1][5] , \stage_1_retimer[1][4] ,
         \stage_1_retimer[1][3] , \stage_1_retimer[1][2] ,
         \stage_1_retimer[1][1] , \stage_1_retimer[1][0] ,
         \stage_1_retimer[0][19] , \stage_1_retimer[0][18] ,
         \stage_1_retimer[0][17] , \stage_1_retimer[0][16] ,
         \stage_1_retimer[0][15] , \stage_1_retimer[0][14] ,
         \stage_1_retimer[0][13] , \stage_1_retimer[0][12] ,
         \stage_1_retimer[0][11] , \stage_1_retimer[0][10] ,
         \stage_1_retimer[0][9] , \stage_1_retimer[0][8] ,
         \stage_1_retimer[0][7] , \stage_1_retimer[0][6] ,
         \stage_1_retimer[0][5] , \stage_1_retimer[0][4] ,
         \stage_1_retimer[0][3] , \stage_1_retimer[0][2] ,
         \stage_1_retimer[0][1] , \stage_1_retimer[0][0] ,
         \stage_2_output[7][19] , \stage_2_output[7][18] ,
         \stage_2_output[7][17] , \stage_2_output[7][16] ,
         \stage_2_output[7][15] , \stage_2_output[7][14] ,
         \stage_2_output[7][13] , \stage_2_output[7][12] ,
         \stage_2_output[7][11] , \stage_2_output[7][10] ,
         \stage_2_output[7][9] , \stage_2_output[7][8] ,
         \stage_2_output[7][7] , \stage_2_output[7][6] ,
         \stage_2_output[7][5] , \stage_2_output[7][4] ,
         \stage_2_output[7][3] , \stage_2_output[7][2] ,
         \stage_2_output[7][1] , \stage_2_output[7][0] ,
         \stage_2_output[6][19] , \stage_2_output[6][18] ,
         \stage_2_output[6][17] , \stage_2_output[6][16] ,
         \stage_2_output[6][15] , \stage_2_output[6][14] ,
         \stage_2_output[6][13] , \stage_2_output[6][12] ,
         \stage_2_output[6][11] , \stage_2_output[6][10] ,
         \stage_2_output[6][9] , \stage_2_output[6][8] ,
         \stage_2_output[6][7] , \stage_2_output[6][6] ,
         \stage_2_output[6][5] , \stage_2_output[6][4] ,
         \stage_2_output[6][3] , \stage_2_output[6][2] ,
         \stage_2_output[6][1] , \stage_2_output[6][0] ,
         \stage_2_output[5][19] , \stage_2_output[5][18] ,
         \stage_2_output[5][17] , \stage_2_output[5][16] ,
         \stage_2_output[5][15] , \stage_2_output[5][14] ,
         \stage_2_output[5][13] , \stage_2_output[5][12] ,
         \stage_2_output[5][11] , \stage_2_output[5][10] ,
         \stage_2_output[5][9] , \stage_2_output[5][8] ,
         \stage_2_output[5][7] , \stage_2_output[5][6] ,
         \stage_2_output[5][5] , \stage_2_output[5][4] ,
         \stage_2_output[5][3] , \stage_2_output[5][2] ,
         \stage_2_output[5][1] , \stage_2_output[5][0] ,
         \stage_2_output[4][19] , \stage_2_output[4][18] ,
         \stage_2_output[4][17] , \stage_2_output[4][16] ,
         \stage_2_output[4][15] , \stage_2_output[4][14] ,
         \stage_2_output[4][13] , \stage_2_output[4][12] ,
         \stage_2_output[4][11] , \stage_2_output[4][10] ,
         \stage_2_output[4][9] , \stage_2_output[4][8] ,
         \stage_2_output[4][7] , \stage_2_output[4][6] ,
         \stage_2_output[4][5] , \stage_2_output[4][4] ,
         \stage_2_output[4][3] , \stage_2_output[4][2] ,
         \stage_2_output[4][1] , \stage_2_output[4][0] ,
         \stage_2_output[3][19] , \stage_2_output[3][18] ,
         \stage_2_output[3][17] , \stage_2_output[3][16] ,
         \stage_2_output[3][15] , \stage_2_output[3][14] ,
         \stage_2_output[3][13] , \stage_2_output[3][12] ,
         \stage_2_output[3][11] , \stage_2_output[3][10] ,
         \stage_2_output[3][9] , \stage_2_output[3][8] ,
         \stage_2_output[3][7] , \stage_2_output[3][6] ,
         \stage_2_output[3][5] , \stage_2_output[3][4] ,
         \stage_2_output[3][3] , \stage_2_output[3][2] ,
         \stage_2_output[3][1] , \stage_2_output[3][0] ,
         \stage_2_output[2][19] , \stage_2_output[2][18] ,
         \stage_2_output[2][17] , \stage_2_output[2][16] ,
         \stage_2_output[2][15] , \stage_2_output[2][14] ,
         \stage_2_output[2][13] , \stage_2_output[2][12] ,
         \stage_2_output[2][11] , \stage_2_output[2][10] ,
         \stage_2_output[2][9] , \stage_2_output[2][8] ,
         \stage_2_output[2][7] , \stage_2_output[2][6] ,
         \stage_2_output[2][5] , \stage_2_output[2][4] ,
         \stage_2_output[2][3] , \stage_2_output[2][2] ,
         \stage_2_output[2][1] , \stage_2_output[2][0] ,
         \stage_2_output[1][19] , \stage_2_output[1][18] ,
         \stage_2_output[1][17] , \stage_2_output[1][16] ,
         \stage_2_output[1][15] , \stage_2_output[1][14] ,
         \stage_2_output[1][13] , \stage_2_output[1][12] ,
         \stage_2_output[1][11] , \stage_2_output[1][10] ,
         \stage_2_output[1][9] , \stage_2_output[1][8] ,
         \stage_2_output[1][7] , \stage_2_output[1][6] ,
         \stage_2_output[1][5] , \stage_2_output[1][4] ,
         \stage_2_output[1][3] , \stage_2_output[1][2] ,
         \stage_2_output[1][1] , \stage_2_output[1][0] ,
         \stage_2_output[0][19] , \stage_2_output[0][18] ,
         \stage_2_output[0][17] , \stage_2_output[0][16] ,
         \stage_2_output[0][15] , \stage_2_output[0][14] ,
         \stage_2_output[0][13] , \stage_2_output[0][12] ,
         \stage_2_output[0][11] , \stage_2_output[0][10] ,
         \stage_2_output[0][9] , \stage_2_output[0][8] ,
         \stage_2_output[0][7] , \stage_2_output[0][6] ,
         \stage_2_output[0][5] , \stage_2_output[0][4] ,
         \stage_2_output[0][3] , \stage_2_output[0][2] ,
         \stage_2_output[0][1] , \stage_2_output[0][0] ,
         \stage_2_retimer[7][19] , \stage_2_retimer[7][18] ,
         \stage_2_retimer[7][17] , \stage_2_retimer[7][16] ,
         \stage_2_retimer[7][15] , \stage_2_retimer[7][14] ,
         \stage_2_retimer[7][13] , \stage_2_retimer[7][12] ,
         \stage_2_retimer[7][11] , \stage_2_retimer[7][10] ,
         \stage_2_retimer[7][9] , \stage_2_retimer[7][8] ,
         \stage_2_retimer[7][7] , \stage_2_retimer[7][6] ,
         \stage_2_retimer[7][5] , \stage_2_retimer[7][4] ,
         \stage_2_retimer[7][3] , \stage_2_retimer[7][2] ,
         \stage_2_retimer[7][1] , \stage_2_retimer[7][0] ,
         \stage_2_retimer[6][19] , \stage_2_retimer[6][18] ,
         \stage_2_retimer[6][17] , \stage_2_retimer[6][16] ,
         \stage_2_retimer[6][15] , \stage_2_retimer[6][14] ,
         \stage_2_retimer[6][13] , \stage_2_retimer[6][12] ,
         \stage_2_retimer[6][11] , \stage_2_retimer[6][10] ,
         \stage_2_retimer[6][9] , \stage_2_retimer[6][8] ,
         \stage_2_retimer[6][7] , \stage_2_retimer[6][6] ,
         \stage_2_retimer[6][5] , \stage_2_retimer[6][4] ,
         \stage_2_retimer[6][3] , \stage_2_retimer[6][2] ,
         \stage_2_retimer[6][1] , \stage_2_retimer[6][0] ,
         \stage_2_retimer[5][19] , \stage_2_retimer[5][18] ,
         \stage_2_retimer[5][17] , \stage_2_retimer[5][16] ,
         \stage_2_retimer[5][15] , \stage_2_retimer[5][14] ,
         \stage_2_retimer[5][13] , \stage_2_retimer[5][12] ,
         \stage_2_retimer[5][11] , \stage_2_retimer[5][10] ,
         \stage_2_retimer[5][9] , \stage_2_retimer[5][8] ,
         \stage_2_retimer[5][7] , \stage_2_retimer[5][6] ,
         \stage_2_retimer[5][5] , \stage_2_retimer[5][4] ,
         \stage_2_retimer[5][3] , \stage_2_retimer[5][2] ,
         \stage_2_retimer[5][1] , \stage_2_retimer[5][0] ,
         \stage_2_retimer[4][19] , \stage_2_retimer[4][18] ,
         \stage_2_retimer[4][17] , \stage_2_retimer[4][16] ,
         \stage_2_retimer[4][15] , \stage_2_retimer[4][14] ,
         \stage_2_retimer[4][13] , \stage_2_retimer[4][12] ,
         \stage_2_retimer[4][11] , \stage_2_retimer[4][10] ,
         \stage_2_retimer[4][9] , \stage_2_retimer[4][8] ,
         \stage_2_retimer[4][7] , \stage_2_retimer[4][6] ,
         \stage_2_retimer[4][5] , \stage_2_retimer[4][4] ,
         \stage_2_retimer[4][3] , \stage_2_retimer[4][2] ,
         \stage_2_retimer[4][1] , \stage_2_retimer[4][0] ,
         \stage_2_retimer[3][19] , \stage_2_retimer[3][18] ,
         \stage_2_retimer[3][17] , \stage_2_retimer[3][16] ,
         \stage_2_retimer[3][15] , \stage_2_retimer[3][14] ,
         \stage_2_retimer[3][13] , \stage_2_retimer[3][12] ,
         \stage_2_retimer[3][11] , \stage_2_retimer[3][10] ,
         \stage_2_retimer[3][9] , \stage_2_retimer[3][8] ,
         \stage_2_retimer[3][7] , \stage_2_retimer[3][6] ,
         \stage_2_retimer[3][5] , \stage_2_retimer[3][4] ,
         \stage_2_retimer[3][3] , \stage_2_retimer[3][2] ,
         \stage_2_retimer[3][1] , \stage_2_retimer[3][0] ,
         \stage_2_retimer[2][19] , \stage_2_retimer[2][18] ,
         \stage_2_retimer[2][17] , \stage_2_retimer[2][16] ,
         \stage_2_retimer[2][15] , \stage_2_retimer[2][14] ,
         \stage_2_retimer[2][13] , \stage_2_retimer[2][12] ,
         \stage_2_retimer[2][11] , \stage_2_retimer[2][10] ,
         \stage_2_retimer[2][9] , \stage_2_retimer[2][8] ,
         \stage_2_retimer[2][7] , \stage_2_retimer[2][6] ,
         \stage_2_retimer[2][5] , \stage_2_retimer[2][4] ,
         \stage_2_retimer[2][3] , \stage_2_retimer[2][2] ,
         \stage_2_retimer[2][1] , \stage_2_retimer[2][0] ,
         \stage_2_retimer[1][19] , \stage_2_retimer[1][18] ,
         \stage_2_retimer[1][17] , \stage_2_retimer[1][16] ,
         \stage_2_retimer[1][15] , \stage_2_retimer[1][14] ,
         \stage_2_retimer[1][13] , \stage_2_retimer[1][12] ,
         \stage_2_retimer[1][11] , \stage_2_retimer[1][10] ,
         \stage_2_retimer[1][9] , \stage_2_retimer[1][8] ,
         \stage_2_retimer[1][7] , \stage_2_retimer[1][6] ,
         \stage_2_retimer[1][5] , \stage_2_retimer[1][4] ,
         \stage_2_retimer[1][3] , \stage_2_retimer[1][2] ,
         \stage_2_retimer[1][1] , \stage_2_retimer[1][0] ,
         \stage_2_retimer[0][19] , \stage_2_retimer[0][18] ,
         \stage_2_retimer[0][17] , \stage_2_retimer[0][16] ,
         \stage_2_retimer[0][15] , \stage_2_retimer[0][14] ,
         \stage_2_retimer[0][13] , \stage_2_retimer[0][12] ,
         \stage_2_retimer[0][11] , \stage_2_retimer[0][10] ,
         \stage_2_retimer[0][9] , \stage_2_retimer[0][8] ,
         \stage_2_retimer[0][7] , \stage_2_retimer[0][6] ,
         \stage_2_retimer[0][5] , \stage_2_retimer[0][4] ,
         \stage_2_retimer[0][3] , \stage_2_retimer[0][2] ,
         \stage_2_retimer[0][1] , \stage_2_retimer[0][0] ,
         \stage_3_output[7][19] , \stage_3_output[7][18] ,
         \stage_3_output[7][17] , \stage_3_output[7][16] ,
         \stage_3_output[7][15] , \stage_3_output[7][14] ,
         \stage_3_output[7][13] , \stage_3_output[7][12] ,
         \stage_3_output[7][11] , \stage_3_output[7][10] ,
         \stage_3_output[7][9] , \stage_3_output[7][8] ,
         \stage_3_output[7][7] , \stage_3_output[7][6] ,
         \stage_3_output[7][5] , \stage_3_output[7][4] ,
         \stage_3_output[7][3] , \stage_3_output[7][2] ,
         \stage_3_output[7][1] , \stage_3_output[7][0] ,
         \stage_3_output[6][19] , \stage_3_output[6][18] ,
         \stage_3_output[6][17] , \stage_3_output[6][16] ,
         \stage_3_output[6][15] , \stage_3_output[6][14] ,
         \stage_3_output[6][13] , \stage_3_output[6][12] ,
         \stage_3_output[6][11] , \stage_3_output[6][10] ,
         \stage_3_output[6][9] , \stage_3_output[6][8] ,
         \stage_3_output[6][7] , \stage_3_output[6][6] ,
         \stage_3_output[6][5] , \stage_3_output[6][4] ,
         \stage_3_output[6][3] , \stage_3_output[6][2] ,
         \stage_3_output[6][1] , \stage_3_output[6][0] ,
         \stage_3_output[5][19] , \stage_3_output[5][18] ,
         \stage_3_output[5][17] , \stage_3_output[5][16] ,
         \stage_3_output[5][15] , \stage_3_output[5][14] ,
         \stage_3_output[5][13] , \stage_3_output[5][12] ,
         \stage_3_output[5][11] , \stage_3_output[5][10] ,
         \stage_3_output[5][9] , \stage_3_output[5][8] ,
         \stage_3_output[5][7] , \stage_3_output[5][6] ,
         \stage_3_output[5][5] , \stage_3_output[5][4] ,
         \stage_3_output[5][3] , \stage_3_output[5][2] ,
         \stage_3_output[5][1] , \stage_3_output[5][0] ,
         \stage_3_output[4][19] , \stage_3_output[4][18] ,
         \stage_3_output[4][17] , \stage_3_output[4][16] ,
         \stage_3_output[4][15] , \stage_3_output[4][14] ,
         \stage_3_output[4][13] , \stage_3_output[4][12] ,
         \stage_3_output[4][11] , \stage_3_output[4][10] ,
         \stage_3_output[4][9] , \stage_3_output[4][8] ,
         \stage_3_output[4][7] , \stage_3_output[4][6] ,
         \stage_3_output[4][5] , \stage_3_output[4][4] ,
         \stage_3_output[4][3] , \stage_3_output[4][2] ,
         \stage_3_output[4][1] , \stage_3_output[4][0] ,
         \stage_3_output[3][19] , \stage_3_output[3][18] ,
         \stage_3_output[3][17] , \stage_3_output[3][16] ,
         \stage_3_output[3][15] , \stage_3_output[3][14] ,
         \stage_3_output[3][13] , \stage_3_output[3][12] ,
         \stage_3_output[3][11] , \stage_3_output[3][10] ,
         \stage_3_output[3][9] , \stage_3_output[3][8] ,
         \stage_3_output[3][7] , \stage_3_output[3][6] ,
         \stage_3_output[3][5] , \stage_3_output[3][4] ,
         \stage_3_output[3][3] , \stage_3_output[3][2] ,
         \stage_3_output[3][1] , \stage_3_output[3][0] ,
         \stage_3_output[2][19] , \stage_3_output[2][18] ,
         \stage_3_output[2][17] , \stage_3_output[2][16] ,
         \stage_3_output[2][15] , \stage_3_output[2][14] ,
         \stage_3_output[2][13] , \stage_3_output[2][12] ,
         \stage_3_output[2][11] , \stage_3_output[2][10] ,
         \stage_3_output[2][9] , \stage_3_output[2][8] ,
         \stage_3_output[2][7] , \stage_3_output[2][6] ,
         \stage_3_output[2][5] , \stage_3_output[2][4] ,
         \stage_3_output[2][3] , \stage_3_output[2][2] ,
         \stage_3_output[2][1] , \stage_3_output[2][0] ,
         \stage_3_output[1][19] , \stage_3_output[1][18] ,
         \stage_3_output[1][17] , \stage_3_output[1][16] ,
         \stage_3_output[1][15] , \stage_3_output[1][14] ,
         \stage_3_output[1][13] , \stage_3_output[1][12] ,
         \stage_3_output[1][11] , \stage_3_output[1][10] ,
         \stage_3_output[1][9] , \stage_3_output[1][8] ,
         \stage_3_output[1][7] , \stage_3_output[1][6] ,
         \stage_3_output[1][5] , \stage_3_output[1][4] ,
         \stage_3_output[1][3] , \stage_3_output[1][2] ,
         \stage_3_output[1][1] , \stage_3_output[1][0] ,
         \stage_3_output[0][19] , \stage_3_output[0][18] ,
         \stage_3_output[0][17] , \stage_3_output[0][16] ,
         \stage_3_output[0][15] , \stage_3_output[0][14] ,
         \stage_3_output[0][13] , \stage_3_output[0][12] ,
         \stage_3_output[0][11] , \stage_3_output[0][10] ,
         \stage_3_output[0][9] , \stage_3_output[0][8] ,
         \stage_3_output[0][7] , \stage_3_output[0][6] ,
         \stage_3_output[0][5] , \stage_3_output[0][4] ,
         \stage_3_output[0][3] , \stage_3_output[0][2] ,
         \stage_3_output[0][1] , \stage_3_output[0][0] ,
         \stage_3_retimer[7][19] , \stage_3_retimer[7][18] ,
         \stage_3_retimer[7][17] , \stage_3_retimer[7][16] ,
         \stage_3_retimer[7][15] , \stage_3_retimer[7][14] ,
         \stage_3_retimer[7][13] , \stage_3_retimer[7][12] ,
         \stage_3_retimer[7][11] , \stage_3_retimer[7][10] ,
         \stage_3_retimer[7][9] , \stage_3_retimer[7][8] ,
         \stage_3_retimer[7][7] , \stage_3_retimer[7][6] ,
         \stage_3_retimer[7][5] , \stage_3_retimer[7][4] ,
         \stage_3_retimer[7][3] , \stage_3_retimer[7][2] ,
         \stage_3_retimer[7][1] , \stage_3_retimer[7][0] ,
         \stage_3_retimer[6][19] , \stage_3_retimer[6][18] ,
         \stage_3_retimer[6][17] , \stage_3_retimer[6][16] ,
         \stage_3_retimer[6][15] , \stage_3_retimer[6][14] ,
         \stage_3_retimer[6][13] , \stage_3_retimer[6][12] ,
         \stage_3_retimer[6][11] , \stage_3_retimer[6][10] ,
         \stage_3_retimer[6][9] , \stage_3_retimer[6][8] ,
         \stage_3_retimer[6][7] , \stage_3_retimer[6][6] ,
         \stage_3_retimer[6][5] , \stage_3_retimer[6][4] ,
         \stage_3_retimer[6][3] , \stage_3_retimer[6][2] ,
         \stage_3_retimer[6][1] , \stage_3_retimer[6][0] ,
         \stage_3_retimer[5][19] , \stage_3_retimer[5][18] ,
         \stage_3_retimer[5][17] , \stage_3_retimer[5][16] ,
         \stage_3_retimer[5][15] , \stage_3_retimer[5][14] ,
         \stage_3_retimer[5][13] , \stage_3_retimer[5][12] ,
         \stage_3_retimer[5][11] , \stage_3_retimer[5][10] ,
         \stage_3_retimer[5][9] , \stage_3_retimer[5][8] ,
         \stage_3_retimer[5][7] , \stage_3_retimer[5][6] ,
         \stage_3_retimer[5][5] , \stage_3_retimer[5][4] ,
         \stage_3_retimer[5][3] , \stage_3_retimer[5][2] ,
         \stage_3_retimer[5][1] , \stage_3_retimer[5][0] ,
         \stage_3_retimer[4][19] , \stage_3_retimer[4][18] ,
         \stage_3_retimer[4][17] , \stage_3_retimer[4][16] ,
         \stage_3_retimer[4][15] , \stage_3_retimer[4][14] ,
         \stage_3_retimer[4][13] , \stage_3_retimer[4][12] ,
         \stage_3_retimer[4][11] , \stage_3_retimer[4][10] ,
         \stage_3_retimer[4][9] , \stage_3_retimer[4][8] ,
         \stage_3_retimer[4][7] , \stage_3_retimer[4][6] ,
         \stage_3_retimer[4][5] , \stage_3_retimer[4][4] ,
         \stage_3_retimer[4][3] , \stage_3_retimer[4][2] ,
         \stage_3_retimer[4][1] , \stage_3_retimer[4][0] ,
         \stage_3_retimer[3][19] , \stage_3_retimer[3][18] ,
         \stage_3_retimer[3][17] , \stage_3_retimer[3][16] ,
         \stage_3_retimer[3][15] , \stage_3_retimer[3][14] ,
         \stage_3_retimer[3][13] , \stage_3_retimer[3][12] ,
         \stage_3_retimer[3][11] , \stage_3_retimer[3][10] ,
         \stage_3_retimer[3][9] , \stage_3_retimer[3][8] ,
         \stage_3_retimer[3][7] , \stage_3_retimer[3][6] ,
         \stage_3_retimer[3][5] , \stage_3_retimer[3][4] ,
         \stage_3_retimer[3][3] , \stage_3_retimer[3][2] ,
         \stage_3_retimer[3][1] , \stage_3_retimer[3][0] ,
         \stage_3_retimer[2][19] , \stage_3_retimer[2][18] ,
         \stage_3_retimer[2][17] , \stage_3_retimer[2][16] ,
         \stage_3_retimer[2][15] , \stage_3_retimer[2][14] ,
         \stage_3_retimer[2][13] , \stage_3_retimer[2][12] ,
         \stage_3_retimer[2][11] , \stage_3_retimer[2][10] ,
         \stage_3_retimer[2][9] , \stage_3_retimer[2][8] ,
         \stage_3_retimer[2][7] , \stage_3_retimer[2][6] ,
         \stage_3_retimer[2][5] , \stage_3_retimer[2][4] ,
         \stage_3_retimer[2][3] , \stage_3_retimer[2][2] ,
         \stage_3_retimer[2][1] , \stage_3_retimer[2][0] ,
         \stage_3_retimer[1][19] , \stage_3_retimer[1][18] ,
         \stage_3_retimer[1][17] , \stage_3_retimer[1][16] ,
         \stage_3_retimer[1][15] , \stage_3_retimer[1][14] ,
         \stage_3_retimer[1][13] , \stage_3_retimer[1][12] ,
         \stage_3_retimer[1][11] , \stage_3_retimer[1][10] ,
         \stage_3_retimer[1][9] , \stage_3_retimer[1][8] ,
         \stage_3_retimer[1][7] , \stage_3_retimer[1][6] ,
         \stage_3_retimer[1][5] , \stage_3_retimer[1][4] ,
         \stage_3_retimer[1][3] , \stage_3_retimer[1][2] ,
         \stage_3_retimer[1][1] , \stage_3_retimer[1][0] ,
         \stage_3_retimer[0][19] , \stage_3_retimer[0][18] ,
         \stage_3_retimer[0][17] , \stage_3_retimer[0][16] ,
         \stage_3_retimer[0][15] , \stage_3_retimer[0][14] ,
         \stage_3_retimer[0][13] , \stage_3_retimer[0][12] ,
         \stage_3_retimer[0][11] , \stage_3_retimer[0][10] ,
         \stage_3_retimer[0][9] , \stage_3_retimer[0][8] ,
         \stage_3_retimer[0][7] , \stage_3_retimer[0][6] ,
         \stage_3_retimer[0][5] , \stage_3_retimer[0][4] ,
         \stage_3_retimer[0][3] , \stage_3_retimer[0][2] ,
         \stage_3_retimer[0][1] , \stage_3_retimer[0][0] ,
         \stage_4_output[7][19] , \stage_4_output[7][18] ,
         \stage_4_output[7][17] , \stage_4_output[7][16] ,
         \stage_4_output[7][15] , \stage_4_output[7][14] ,
         \stage_4_output[7][13] , \stage_4_output[7][12] ,
         \stage_4_output[7][11] , \stage_4_output[7][10] ,
         \stage_4_output[7][9] , \stage_4_output[7][8] ,
         \stage_4_output[7][7] , \stage_4_output[7][6] ,
         \stage_4_output[7][5] , \stage_4_output[7][4] ,
         \stage_4_output[7][3] , \stage_4_output[7][2] ,
         \stage_4_output[7][1] , \stage_4_output[7][0] ,
         \stage_4_output[6][19] , \stage_4_output[6][18] ,
         \stage_4_output[6][17] , \stage_4_output[6][16] ,
         \stage_4_output[6][15] , \stage_4_output[6][14] ,
         \stage_4_output[6][13] , \stage_4_output[6][12] ,
         \stage_4_output[6][11] , \stage_4_output[6][10] ,
         \stage_4_output[6][9] , \stage_4_output[6][8] ,
         \stage_4_output[6][7] , \stage_4_output[6][6] ,
         \stage_4_output[6][5] , \stage_4_output[6][4] ,
         \stage_4_output[6][3] , \stage_4_output[6][2] ,
         \stage_4_output[6][1] , \stage_4_output[6][0] ,
         \stage_4_output[5][19] , \stage_4_output[5][18] ,
         \stage_4_output[5][17] , \stage_4_output[5][16] ,
         \stage_4_output[5][15] , \stage_4_output[5][14] ,
         \stage_4_output[5][13] , \stage_4_output[5][12] ,
         \stage_4_output[5][11] , \stage_4_output[5][10] ,
         \stage_4_output[5][9] , \stage_4_output[5][8] ,
         \stage_4_output[5][7] , \stage_4_output[5][6] ,
         \stage_4_output[5][5] , \stage_4_output[5][4] ,
         \stage_4_output[5][3] , \stage_4_output[5][2] ,
         \stage_4_output[5][1] , \stage_4_output[5][0] ,
         \stage_4_output[4][19] , \stage_4_output[4][18] ,
         \stage_4_output[4][17] , \stage_4_output[4][16] ,
         \stage_4_output[4][15] , \stage_4_output[4][14] ,
         \stage_4_output[4][13] , \stage_4_output[4][12] ,
         \stage_4_output[4][11] , \stage_4_output[4][10] ,
         \stage_4_output[4][9] , \stage_4_output[4][8] ,
         \stage_4_output[4][7] , \stage_4_output[4][6] ,
         \stage_4_output[4][5] , \stage_4_output[4][4] ,
         \stage_4_output[4][3] , \stage_4_output[4][2] ,
         \stage_4_output[4][1] , \stage_4_output[4][0] ,
         \stage_4_output[3][19] , \stage_4_output[3][18] ,
         \stage_4_output[3][17] , \stage_4_output[3][16] ,
         \stage_4_output[3][15] , \stage_4_output[3][14] ,
         \stage_4_output[3][13] , \stage_4_output[3][12] ,
         \stage_4_output[3][11] , \stage_4_output[3][10] ,
         \stage_4_output[3][9] , \stage_4_output[3][8] ,
         \stage_4_output[3][7] , \stage_4_output[3][6] ,
         \stage_4_output[3][5] , \stage_4_output[3][4] ,
         \stage_4_output[3][3] , \stage_4_output[3][2] ,
         \stage_4_output[3][1] , \stage_4_output[3][0] ,
         \stage_4_output[2][19] , \stage_4_output[2][18] ,
         \stage_4_output[2][17] , \stage_4_output[2][16] ,
         \stage_4_output[2][15] , \stage_4_output[2][14] ,
         \stage_4_output[2][13] , \stage_4_output[2][12] ,
         \stage_4_output[2][11] , \stage_4_output[2][10] ,
         \stage_4_output[2][9] , \stage_4_output[2][8] ,
         \stage_4_output[2][7] , \stage_4_output[2][6] ,
         \stage_4_output[2][5] , \stage_4_output[2][4] ,
         \stage_4_output[2][3] , \stage_4_output[2][2] ,
         \stage_4_output[2][1] , \stage_4_output[2][0] ,
         \stage_4_output[1][19] , \stage_4_output[1][18] ,
         \stage_4_output[1][17] , \stage_4_output[1][16] ,
         \stage_4_output[1][15] , \stage_4_output[1][14] ,
         \stage_4_output[1][13] , \stage_4_output[1][12] ,
         \stage_4_output[1][11] , \stage_4_output[1][10] ,
         \stage_4_output[1][9] , \stage_4_output[1][8] ,
         \stage_4_output[1][7] , \stage_4_output[1][6] ,
         \stage_4_output[1][5] , \stage_4_output[1][4] ,
         \stage_4_output[1][3] , \stage_4_output[1][2] ,
         \stage_4_output[1][1] , \stage_4_output[1][0] ,
         \stage_4_output[0][19] , \stage_4_output[0][18] ,
         \stage_4_output[0][17] , \stage_4_output[0][16] ,
         \stage_4_output[0][15] , \stage_4_output[0][14] ,
         \stage_4_output[0][13] , \stage_4_output[0][12] ,
         \stage_4_output[0][11] , \stage_4_output[0][10] ,
         \stage_4_output[0][9] , \stage_4_output[0][8] ,
         \stage_4_output[0][7] , \stage_4_output[0][6] ,
         \stage_4_output[0][5] , \stage_4_output[0][4] ,
         \stage_4_output[0][3] , \stage_4_output[0][2] ,
         \stage_4_output[0][1] , \stage_4_output[0][0] ;
  assign \in_upper_00[3]  = port_en_n[0];
  assign \in_lower_00[3]  = port_en_n[1];
  assign \in_upper_01[3]  = port_en_n[2];
  assign \in_lower_01[3]  = port_en_n[3];
  assign in_upper_02_3 = port_en_n[4];
  assign \in_lower_02[3]  = port_en_n[5];
  assign \in_upper_03[3]  = port_en_n[6];

  crossbar_0 u_00_crossbar ( .in_upper({in_input[127:112], \in_upper_00[3] , 
        \in_upper_00[3] , \in_upper_00[3] , \in_upper_00[3] }), .in_lower({
        in_input[111:96], \in_lower_00[3] , \in_lower_00[3] , \in_lower_00[3] , 
        \*Logic1* }), .in_control(in_control[19]), .out_upper({
        \stage_0_output[0][19] , \stage_0_output[0][18] , 
        \stage_0_output[0][17] , \stage_0_output[0][16] , 
        \stage_0_output[0][15] , \stage_0_output[0][14] , 
        \stage_0_output[0][13] , \stage_0_output[0][12] , 
        \stage_0_output[0][11] , \stage_0_output[0][10] , 
        \stage_0_output[0][9] , \stage_0_output[0][8] , \stage_0_output[0][7] , 
        \stage_0_output[0][6] , \stage_0_output[0][5] , \stage_0_output[0][4] , 
        \stage_0_output[0][3] , \stage_0_output[0][2] , \stage_0_output[0][1] , 
        \stage_0_output[0][0] }), .out_lower({\stage_0_output[1][19] , 
        \stage_0_output[1][18] , \stage_0_output[1][17] , 
        \stage_0_output[1][16] , \stage_0_output[1][15] , 
        \stage_0_output[1][14] , \stage_0_output[1][13] , 
        \stage_0_output[1][12] , \stage_0_output[1][11] , 
        \stage_0_output[1][10] , \stage_0_output[1][9] , 
        \stage_0_output[1][8] , \stage_0_output[1][7] , \stage_0_output[1][6] , 
        \stage_0_output[1][5] , \stage_0_output[1][4] , \stage_0_output[1][3] , 
        \stage_0_output[1][2] , \stage_0_output[1][1] , \stage_0_output[1][0] }) );
  crossbar_19 u_01_crossbar ( .in_upper({in_input[95:80], \in_upper_01[3] , 
        \in_upper_01[3] , \*Logic1* , \in_upper_01[3] }), .in_lower({
        in_input[79:64], \in_lower_01[3] , \in_lower_01[3] , \*Logic1* , 
        \*Logic1* }), .in_control(in_control[18]), .out_upper({
        \stage_0_output[2][19] , \stage_0_output[2][18] , 
        \stage_0_output[2][17] , \stage_0_output[2][16] , 
        \stage_0_output[2][15] , \stage_0_output[2][14] , 
        \stage_0_output[2][13] , \stage_0_output[2][12] , 
        \stage_0_output[2][11] , \stage_0_output[2][10] , 
        \stage_0_output[2][9] , \stage_0_output[2][8] , \stage_0_output[2][7] , 
        \stage_0_output[2][6] , \stage_0_output[2][5] , \stage_0_output[2][4] , 
        \stage_0_output[2][3] , \stage_0_output[2][2] , \stage_0_output[2][1] , 
        \stage_0_output[2][0] }), .out_lower({\stage_0_output[3][19] , 
        \stage_0_output[3][18] , \stage_0_output[3][17] , 
        \stage_0_output[3][16] , \stage_0_output[3][15] , 
        \stage_0_output[3][14] , \stage_0_output[3][13] , 
        \stage_0_output[3][12] , \stage_0_output[3][11] , 
        \stage_0_output[3][10] , \stage_0_output[3][9] , 
        \stage_0_output[3][8] , \stage_0_output[3][7] , \stage_0_output[3][6] , 
        \stage_0_output[3][5] , \stage_0_output[3][4] , \stage_0_output[3][3] , 
        \stage_0_output[3][2] , \stage_0_output[3][1] , \stage_0_output[3][0] }) );
  crossbar_18 u_02_crossbar ( .in_upper({in_input[63:48], in_upper_02_3, 
        \*Logic1* , in_upper_02_3, in_upper_02_3}), .in_lower({in_input[47:32], 
        \in_lower_02[3] , \*Logic1* , \in_lower_02[3] , \*Logic1* }), 
        .in_control(in_control[17]), .out_upper({\stage_0_output[4][19] , 
        \stage_0_output[4][18] , \stage_0_output[4][17] , 
        \stage_0_output[4][16] , \stage_0_output[4][15] , 
        \stage_0_output[4][14] , \stage_0_output[4][13] , 
        \stage_0_output[4][12] , \stage_0_output[4][11] , 
        \stage_0_output[4][10] , \stage_0_output[4][9] , 
        \stage_0_output[4][8] , \stage_0_output[4][7] , \stage_0_output[4][6] , 
        \stage_0_output[4][5] , \stage_0_output[4][4] , \stage_0_output[4][3] , 
        \stage_0_output[4][2] , \stage_0_output[4][1] , \stage_0_output[4][0] }), .out_lower({\stage_0_output[5][19] , \stage_0_output[5][18] , 
        \stage_0_output[5][17] , \stage_0_output[5][16] , 
        \stage_0_output[5][15] , \stage_0_output[5][14] , 
        \stage_0_output[5][13] , \stage_0_output[5][12] , 
        \stage_0_output[5][11] , \stage_0_output[5][10] , 
        \stage_0_output[5][9] , \stage_0_output[5][8] , \stage_0_output[5][7] , 
        \stage_0_output[5][6] , \stage_0_output[5][5] , \stage_0_output[5][4] , 
        \stage_0_output[5][3] , \stage_0_output[5][2] , \stage_0_output[5][1] , 
        \stage_0_output[5][0] }) );
  crossbar_17 u_03_crossbar ( .in_upper({in_input[31:16], \in_upper_03[3] , 
        \*Logic1* , \*Logic1* , \in_upper_03[3] }), .in_lower({in_input[15:0], 
        port_en_n[7], \*Logic1* , \*Logic1* , \*Logic1* }), .in_control(
        in_control[16]), .out_upper({\stage_0_output[6][19] , 
        \stage_0_output[6][18] , \stage_0_output[6][17] , 
        \stage_0_output[6][16] , \stage_0_output[6][15] , 
        \stage_0_output[6][14] , \stage_0_output[6][13] , 
        \stage_0_output[6][12] , \stage_0_output[6][11] , 
        \stage_0_output[6][10] , \stage_0_output[6][9] , 
        \stage_0_output[6][8] , \stage_0_output[6][7] , \stage_0_output[6][6] , 
        \stage_0_output[6][5] , \stage_0_output[6][4] , \stage_0_output[6][3] , 
        \stage_0_output[6][2] , \stage_0_output[6][1] , \stage_0_output[6][0] }), .out_lower({\stage_0_output[7][19] , \stage_0_output[7][18] , 
        \stage_0_output[7][17] , \stage_0_output[7][16] , 
        \stage_0_output[7][15] , \stage_0_output[7][14] , 
        \stage_0_output[7][13] , \stage_0_output[7][12] , 
        \stage_0_output[7][11] , \stage_0_output[7][10] , 
        \stage_0_output[7][9] , \stage_0_output[7][8] , \stage_0_output[7][7] , 
        \stage_0_output[7][6] , \stage_0_output[7][5] , \stage_0_output[7][4] , 
        \stage_0_output[7][3] , \stage_0_output[7][2] , \stage_0_output[7][1] , 
        \stage_0_output[7][0] }) );
  crossbar_16 u_10_crossbar ( .in_upper({\stage_0_retimer[0][19] , 
        \stage_0_retimer[0][18] , \stage_0_retimer[0][17] , 
        \stage_0_retimer[0][16] , \stage_0_retimer[0][15] , 
        \stage_0_retimer[0][14] , \stage_0_retimer[0][13] , 
        \stage_0_retimer[0][12] , \stage_0_retimer[0][11] , 
        \stage_0_retimer[0][10] , \stage_0_retimer[0][9] , 
        \stage_0_retimer[0][8] , \stage_0_retimer[0][7] , 
        \stage_0_retimer[0][6] , \stage_0_retimer[0][5] , 
        \stage_0_retimer[0][4] , \stage_0_retimer[0][3] , 
        \stage_0_retimer[0][2] , \stage_0_retimer[0][1] , 
        \stage_0_retimer[0][0] }), .in_lower({\stage_0_retimer[2][19] , 
        \stage_0_retimer[2][18] , \stage_0_retimer[2][17] , 
        \stage_0_retimer[2][16] , \stage_0_retimer[2][15] , 
        \stage_0_retimer[2][14] , \stage_0_retimer[2][13] , 
        \stage_0_retimer[2][12] , \stage_0_retimer[2][11] , 
        \stage_0_retimer[2][10] , \stage_0_retimer[2][9] , 
        \stage_0_retimer[2][8] , \stage_0_retimer[2][7] , 
        \stage_0_retimer[2][6] , \stage_0_retimer[2][5] , 
        \stage_0_retimer[2][4] , \stage_0_retimer[2][3] , 
        \stage_0_retimer[2][2] , \stage_0_retimer[2][1] , 
        \stage_0_retimer[2][0] }), .in_control(in_control[15]), .out_upper({
        \stage_1_output[0][19] , \stage_1_output[0][18] , 
        \stage_1_output[0][17] , \stage_1_output[0][16] , 
        \stage_1_output[0][15] , \stage_1_output[0][14] , 
        \stage_1_output[0][13] , \stage_1_output[0][12] , 
        \stage_1_output[0][11] , \stage_1_output[0][10] , 
        \stage_1_output[0][9] , \stage_1_output[0][8] , \stage_1_output[0][7] , 
        \stage_1_output[0][6] , \stage_1_output[0][5] , \stage_1_output[0][4] , 
        \stage_1_output[0][3] , \stage_1_output[0][2] , \stage_1_output[0][1] , 
        \stage_1_output[0][0] }), .out_lower({\stage_1_output[1][19] , 
        \stage_1_output[1][18] , \stage_1_output[1][17] , 
        \stage_1_output[1][16] , \stage_1_output[1][15] , 
        \stage_1_output[1][14] , \stage_1_output[1][13] , 
        \stage_1_output[1][12] , \stage_1_output[1][11] , 
        \stage_1_output[1][10] , \stage_1_output[1][9] , 
        \stage_1_output[1][8] , \stage_1_output[1][7] , \stage_1_output[1][6] , 
        \stage_1_output[1][5] , \stage_1_output[1][4] , \stage_1_output[1][3] , 
        \stage_1_output[1][2] , \stage_1_output[1][1] , \stage_1_output[1][0] }) );
  crossbar_15 u_11_crossbar ( .in_upper({\stage_0_retimer[4][19] , 
        \stage_0_retimer[4][18] , \stage_0_retimer[4][17] , 
        \stage_0_retimer[4][16] , \stage_0_retimer[4][15] , 
        \stage_0_retimer[4][14] , \stage_0_retimer[4][13] , 
        \stage_0_retimer[4][12] , \stage_0_retimer[4][11] , 
        \stage_0_retimer[4][10] , \stage_0_retimer[4][9] , 
        \stage_0_retimer[4][8] , \stage_0_retimer[4][7] , 
        \stage_0_retimer[4][6] , \stage_0_retimer[4][5] , 
        \stage_0_retimer[4][4] , \stage_0_retimer[4][3] , 
        \stage_0_retimer[4][2] , \stage_0_retimer[4][1] , 
        \stage_0_retimer[4][0] }), .in_lower({\stage_0_retimer[6][19] , 
        \stage_0_retimer[6][18] , \stage_0_retimer[6][17] , 
        \stage_0_retimer[6][16] , \stage_0_retimer[6][15] , 
        \stage_0_retimer[6][14] , \stage_0_retimer[6][13] , 
        \stage_0_retimer[6][12] , \stage_0_retimer[6][11] , 
        \stage_0_retimer[6][10] , \stage_0_retimer[6][9] , 
        \stage_0_retimer[6][8] , \stage_0_retimer[6][7] , 
        \stage_0_retimer[6][6] , \stage_0_retimer[6][5] , 
        \stage_0_retimer[6][4] , \stage_0_retimer[6][3] , 
        \stage_0_retimer[6][2] , \stage_0_retimer[6][1] , 
        \stage_0_retimer[6][0] }), .in_control(in_control[14]), .out_upper({
        \stage_1_output[2][19] , \stage_1_output[2][18] , 
        \stage_1_output[2][17] , \stage_1_output[2][16] , 
        \stage_1_output[2][15] , \stage_1_output[2][14] , 
        \stage_1_output[2][13] , \stage_1_output[2][12] , 
        \stage_1_output[2][11] , \stage_1_output[2][10] , 
        \stage_1_output[2][9] , \stage_1_output[2][8] , \stage_1_output[2][7] , 
        \stage_1_output[2][6] , \stage_1_output[2][5] , \stage_1_output[2][4] , 
        \stage_1_output[2][3] , \stage_1_output[2][2] , \stage_1_output[2][1] , 
        \stage_1_output[2][0] }), .out_lower({\stage_1_output[3][19] , 
        \stage_1_output[3][18] , \stage_1_output[3][17] , 
        \stage_1_output[3][16] , \stage_1_output[3][15] , 
        \stage_1_output[3][14] , \stage_1_output[3][13] , 
        \stage_1_output[3][12] , \stage_1_output[3][11] , 
        \stage_1_output[3][10] , \stage_1_output[3][9] , 
        \stage_1_output[3][8] , \stage_1_output[3][7] , \stage_1_output[3][6] , 
        \stage_1_output[3][5] , \stage_1_output[3][4] , \stage_1_output[3][3] , 
        \stage_1_output[3][2] , \stage_1_output[3][1] , \stage_1_output[3][0] }) );
  crossbar_14 u_12_crossbar ( .in_upper({\stage_0_retimer[1][19] , 
        \stage_0_retimer[1][18] , \stage_0_retimer[1][17] , 
        \stage_0_retimer[1][16] , \stage_0_retimer[1][15] , 
        \stage_0_retimer[1][14] , \stage_0_retimer[1][13] , 
        \stage_0_retimer[1][12] , \stage_0_retimer[1][11] , 
        \stage_0_retimer[1][10] , \stage_0_retimer[1][9] , 
        \stage_0_retimer[1][8] , \stage_0_retimer[1][7] , 
        \stage_0_retimer[1][6] , \stage_0_retimer[1][5] , 
        \stage_0_retimer[1][4] , \stage_0_retimer[1][3] , 
        \stage_0_retimer[1][2] , \stage_0_retimer[1][1] , 
        \stage_0_retimer[1][0] }), .in_lower({\stage_0_retimer[3][19] , 
        \stage_0_retimer[3][18] , \stage_0_retimer[3][17] , 
        \stage_0_retimer[3][16] , \stage_0_retimer[3][15] , 
        \stage_0_retimer[3][14] , \stage_0_retimer[3][13] , 
        \stage_0_retimer[3][12] , \stage_0_retimer[3][11] , 
        \stage_0_retimer[3][10] , \stage_0_retimer[3][9] , 
        \stage_0_retimer[3][8] , \stage_0_retimer[3][7] , 
        \stage_0_retimer[3][6] , \stage_0_retimer[3][5] , 
        \stage_0_retimer[3][4] , \stage_0_retimer[3][3] , 
        \stage_0_retimer[3][2] , \stage_0_retimer[3][1] , 
        \stage_0_retimer[3][0] }), .in_control(in_control[13]), .out_upper({
        \stage_1_output[4][19] , \stage_1_output[4][18] , 
        \stage_1_output[4][17] , \stage_1_output[4][16] , 
        \stage_1_output[4][15] , \stage_1_output[4][14] , 
        \stage_1_output[4][13] , \stage_1_output[4][12] , 
        \stage_1_output[4][11] , \stage_1_output[4][10] , 
        \stage_1_output[4][9] , \stage_1_output[4][8] , \stage_1_output[4][7] , 
        \stage_1_output[4][6] , \stage_1_output[4][5] , \stage_1_output[4][4] , 
        \stage_1_output[4][3] , \stage_1_output[4][2] , \stage_1_output[4][1] , 
        \stage_1_output[4][0] }), .out_lower({\stage_1_output[5][19] , 
        \stage_1_output[5][18] , \stage_1_output[5][17] , 
        \stage_1_output[5][16] , \stage_1_output[5][15] , 
        \stage_1_output[5][14] , \stage_1_output[5][13] , 
        \stage_1_output[5][12] , \stage_1_output[5][11] , 
        \stage_1_output[5][10] , \stage_1_output[5][9] , 
        \stage_1_output[5][8] , \stage_1_output[5][7] , \stage_1_output[5][6] , 
        \stage_1_output[5][5] , \stage_1_output[5][4] , \stage_1_output[5][3] , 
        \stage_1_output[5][2] , \stage_1_output[5][1] , \stage_1_output[5][0] }) );
  crossbar_13 u_13_crossbar ( .in_upper({\stage_0_retimer[5][19] , 
        \stage_0_retimer[5][18] , \stage_0_retimer[5][17] , 
        \stage_0_retimer[5][16] , \stage_0_retimer[5][15] , 
        \stage_0_retimer[5][14] , \stage_0_retimer[5][13] , 
        \stage_0_retimer[5][12] , \stage_0_retimer[5][11] , 
        \stage_0_retimer[5][10] , \stage_0_retimer[5][9] , 
        \stage_0_retimer[5][8] , \stage_0_retimer[5][7] , 
        \stage_0_retimer[5][6] , \stage_0_retimer[5][5] , 
        \stage_0_retimer[5][4] , \stage_0_retimer[5][3] , 
        \stage_0_retimer[5][2] , \stage_0_retimer[5][1] , 
        \stage_0_retimer[5][0] }), .in_lower({\stage_0_retimer[7][19] , 
        \stage_0_retimer[7][18] , \stage_0_retimer[7][17] , 
        \stage_0_retimer[7][16] , \stage_0_retimer[7][15] , 
        \stage_0_retimer[7][14] , \stage_0_retimer[7][13] , 
        \stage_0_retimer[7][12] , \stage_0_retimer[7][11] , 
        \stage_0_retimer[7][10] , \stage_0_retimer[7][9] , 
        \stage_0_retimer[7][8] , \stage_0_retimer[7][7] , 
        \stage_0_retimer[7][6] , \stage_0_retimer[7][5] , 
        \stage_0_retimer[7][4] , \stage_0_retimer[7][3] , 
        \stage_0_retimer[7][2] , \stage_0_retimer[7][1] , 
        \stage_0_retimer[7][0] }), .in_control(in_control[12]), .out_upper({
        \stage_1_output[6][19] , \stage_1_output[6][18] , 
        \stage_1_output[6][17] , \stage_1_output[6][16] , 
        \stage_1_output[6][15] , \stage_1_output[6][14] , 
        \stage_1_output[6][13] , \stage_1_output[6][12] , 
        \stage_1_output[6][11] , \stage_1_output[6][10] , 
        \stage_1_output[6][9] , \stage_1_output[6][8] , \stage_1_output[6][7] , 
        \stage_1_output[6][6] , \stage_1_output[6][5] , \stage_1_output[6][4] , 
        \stage_1_output[6][3] , \stage_1_output[6][2] , \stage_1_output[6][1] , 
        \stage_1_output[6][0] }), .out_lower({\stage_1_output[7][19] , 
        \stage_1_output[7][18] , \stage_1_output[7][17] , 
        \stage_1_output[7][16] , \stage_1_output[7][15] , 
        \stage_1_output[7][14] , \stage_1_output[7][13] , 
        \stage_1_output[7][12] , \stage_1_output[7][11] , 
        \stage_1_output[7][10] , \stage_1_output[7][9] , 
        \stage_1_output[7][8] , \stage_1_output[7][7] , \stage_1_output[7][6] , 
        \stage_1_output[7][5] , \stage_1_output[7][4] , \stage_1_output[7][3] , 
        \stage_1_output[7][2] , \stage_1_output[7][1] , \stage_1_output[7][0] }) );
  crossbar_12 u_20_crossbar ( .in_upper({\stage_1_retimer[0][19] , 
        \stage_1_retimer[0][18] , \stage_1_retimer[0][17] , 
        \stage_1_retimer[0][16] , \stage_1_retimer[0][15] , 
        \stage_1_retimer[0][14] , \stage_1_retimer[0][13] , 
        \stage_1_retimer[0][12] , \stage_1_retimer[0][11] , 
        \stage_1_retimer[0][10] , \stage_1_retimer[0][9] , 
        \stage_1_retimer[0][8] , \stage_1_retimer[0][7] , 
        \stage_1_retimer[0][6] , \stage_1_retimer[0][5] , 
        \stage_1_retimer[0][4] , \stage_1_retimer[0][3] , 
        \stage_1_retimer[0][2] , \stage_1_retimer[0][1] , 
        \stage_1_retimer[0][0] }), .in_lower({\stage_1_retimer[2][19] , 
        \stage_1_retimer[2][18] , \stage_1_retimer[2][17] , 
        \stage_1_retimer[2][16] , \stage_1_retimer[2][15] , 
        \stage_1_retimer[2][14] , \stage_1_retimer[2][13] , 
        \stage_1_retimer[2][12] , \stage_1_retimer[2][11] , 
        \stage_1_retimer[2][10] , \stage_1_retimer[2][9] , 
        \stage_1_retimer[2][8] , \stage_1_retimer[2][7] , 
        \stage_1_retimer[2][6] , \stage_1_retimer[2][5] , 
        \stage_1_retimer[2][4] , \stage_1_retimer[2][3] , 
        \stage_1_retimer[2][2] , \stage_1_retimer[2][1] , 
        \stage_1_retimer[2][0] }), .in_control(in_control[11]), .out_upper({
        \stage_2_output[0][19] , \stage_2_output[0][18] , 
        \stage_2_output[0][17] , \stage_2_output[0][16] , 
        \stage_2_output[0][15] , \stage_2_output[0][14] , 
        \stage_2_output[0][13] , \stage_2_output[0][12] , 
        \stage_2_output[0][11] , \stage_2_output[0][10] , 
        \stage_2_output[0][9] , \stage_2_output[0][8] , \stage_2_output[0][7] , 
        \stage_2_output[0][6] , \stage_2_output[0][5] , \stage_2_output[0][4] , 
        \stage_2_output[0][3] , \stage_2_output[0][2] , \stage_2_output[0][1] , 
        \stage_2_output[0][0] }), .out_lower({\stage_2_output[1][19] , 
        \stage_2_output[1][18] , \stage_2_output[1][17] , 
        \stage_2_output[1][16] , \stage_2_output[1][15] , 
        \stage_2_output[1][14] , \stage_2_output[1][13] , 
        \stage_2_output[1][12] , \stage_2_output[1][11] , 
        \stage_2_output[1][10] , \stage_2_output[1][9] , 
        \stage_2_output[1][8] , \stage_2_output[1][7] , \stage_2_output[1][6] , 
        \stage_2_output[1][5] , \stage_2_output[1][4] , \stage_2_output[1][3] , 
        \stage_2_output[1][2] , \stage_2_output[1][1] , \stage_2_output[1][0] }) );
  crossbar_11 u_21_crossbar ( .in_upper({\stage_1_retimer[1][19] , 
        \stage_1_retimer[1][18] , \stage_1_retimer[1][17] , 
        \stage_1_retimer[1][16] , \stage_1_retimer[1][15] , 
        \stage_1_retimer[1][14] , \stage_1_retimer[1][13] , 
        \stage_1_retimer[1][12] , \stage_1_retimer[1][11] , 
        \stage_1_retimer[1][10] , \stage_1_retimer[1][9] , 
        \stage_1_retimer[1][8] , \stage_1_retimer[1][7] , 
        \stage_1_retimer[1][6] , \stage_1_retimer[1][5] , 
        \stage_1_retimer[1][4] , \stage_1_retimer[1][3] , 
        \stage_1_retimer[1][2] , \stage_1_retimer[1][1] , 
        \stage_1_retimer[1][0] }), .in_lower({\stage_1_retimer[3][19] , 
        \stage_1_retimer[3][18] , \stage_1_retimer[3][17] , 
        \stage_1_retimer[3][16] , \stage_1_retimer[3][15] , 
        \stage_1_retimer[3][14] , \stage_1_retimer[3][13] , 
        \stage_1_retimer[3][12] , \stage_1_retimer[3][11] , 
        \stage_1_retimer[3][10] , \stage_1_retimer[3][9] , 
        \stage_1_retimer[3][8] , \stage_1_retimer[3][7] , 
        \stage_1_retimer[3][6] , \stage_1_retimer[3][5] , 
        \stage_1_retimer[3][4] , \stage_1_retimer[3][3] , 
        \stage_1_retimer[3][2] , \stage_1_retimer[3][1] , 
        \stage_1_retimer[3][0] }), .in_control(in_control[10]), .out_upper({
        \stage_2_output[2][19] , \stage_2_output[2][18] , 
        \stage_2_output[2][17] , \stage_2_output[2][16] , 
        \stage_2_output[2][15] , \stage_2_output[2][14] , 
        \stage_2_output[2][13] , \stage_2_output[2][12] , 
        \stage_2_output[2][11] , \stage_2_output[2][10] , 
        \stage_2_output[2][9] , \stage_2_output[2][8] , \stage_2_output[2][7] , 
        \stage_2_output[2][6] , \stage_2_output[2][5] , \stage_2_output[2][4] , 
        \stage_2_output[2][3] , \stage_2_output[2][2] , \stage_2_output[2][1] , 
        \stage_2_output[2][0] }), .out_lower({\stage_2_output[3][19] , 
        \stage_2_output[3][18] , \stage_2_output[3][17] , 
        \stage_2_output[3][16] , \stage_2_output[3][15] , 
        \stage_2_output[3][14] , \stage_2_output[3][13] , 
        \stage_2_output[3][12] , \stage_2_output[3][11] , 
        \stage_2_output[3][10] , \stage_2_output[3][9] , 
        \stage_2_output[3][8] , \stage_2_output[3][7] , \stage_2_output[3][6] , 
        \stage_2_output[3][5] , \stage_2_output[3][4] , \stage_2_output[3][3] , 
        \stage_2_output[3][2] , \stage_2_output[3][1] , \stage_2_output[3][0] }) );
  crossbar_10 u_22_crossbar ( .in_upper({\stage_1_retimer[4][19] , 
        \stage_1_retimer[4][18] , \stage_1_retimer[4][17] , 
        \stage_1_retimer[4][16] , \stage_1_retimer[4][15] , 
        \stage_1_retimer[4][14] , \stage_1_retimer[4][13] , 
        \stage_1_retimer[4][12] , \stage_1_retimer[4][11] , 
        \stage_1_retimer[4][10] , \stage_1_retimer[4][9] , 
        \stage_1_retimer[4][8] , \stage_1_retimer[4][7] , 
        \stage_1_retimer[4][6] , \stage_1_retimer[4][5] , 
        \stage_1_retimer[4][4] , \stage_1_retimer[4][3] , 
        \stage_1_retimer[4][2] , \stage_1_retimer[4][1] , 
        \stage_1_retimer[4][0] }), .in_lower({\stage_1_retimer[6][19] , 
        \stage_1_retimer[6][18] , \stage_1_retimer[6][17] , 
        \stage_1_retimer[6][16] , \stage_1_retimer[6][15] , 
        \stage_1_retimer[6][14] , \stage_1_retimer[6][13] , 
        \stage_1_retimer[6][12] , \stage_1_retimer[6][11] , 
        \stage_1_retimer[6][10] , \stage_1_retimer[6][9] , 
        \stage_1_retimer[6][8] , \stage_1_retimer[6][7] , 
        \stage_1_retimer[6][6] , \stage_1_retimer[6][5] , 
        \stage_1_retimer[6][4] , \stage_1_retimer[6][3] , 
        \stage_1_retimer[6][2] , \stage_1_retimer[6][1] , 
        \stage_1_retimer[6][0] }), .in_control(in_control[9]), .out_upper({
        \stage_2_output[4][19] , \stage_2_output[4][18] , 
        \stage_2_output[4][17] , \stage_2_output[4][16] , 
        \stage_2_output[4][15] , \stage_2_output[4][14] , 
        \stage_2_output[4][13] , \stage_2_output[4][12] , 
        \stage_2_output[4][11] , \stage_2_output[4][10] , 
        \stage_2_output[4][9] , \stage_2_output[4][8] , \stage_2_output[4][7] , 
        \stage_2_output[4][6] , \stage_2_output[4][5] , \stage_2_output[4][4] , 
        \stage_2_output[4][3] , \stage_2_output[4][2] , \stage_2_output[4][1] , 
        \stage_2_output[4][0] }), .out_lower({\stage_2_output[5][19] , 
        \stage_2_output[5][18] , \stage_2_output[5][17] , 
        \stage_2_output[5][16] , \stage_2_output[5][15] , 
        \stage_2_output[5][14] , \stage_2_output[5][13] , 
        \stage_2_output[5][12] , \stage_2_output[5][11] , 
        \stage_2_output[5][10] , \stage_2_output[5][9] , 
        \stage_2_output[5][8] , \stage_2_output[5][7] , \stage_2_output[5][6] , 
        \stage_2_output[5][5] , \stage_2_output[5][4] , \stage_2_output[5][3] , 
        \stage_2_output[5][2] , \stage_2_output[5][1] , \stage_2_output[5][0] }) );
  crossbar_9 u_23_crossbar ( .in_upper({\stage_1_retimer[5][19] , 
        \stage_1_retimer[5][18] , \stage_1_retimer[5][17] , 
        \stage_1_retimer[5][16] , \stage_1_retimer[5][15] , 
        \stage_1_retimer[5][14] , \stage_1_retimer[5][13] , 
        \stage_1_retimer[5][12] , \stage_1_retimer[5][11] , 
        \stage_1_retimer[5][10] , \stage_1_retimer[5][9] , 
        \stage_1_retimer[5][8] , \stage_1_retimer[5][7] , 
        \stage_1_retimer[5][6] , \stage_1_retimer[5][5] , 
        \stage_1_retimer[5][4] , \stage_1_retimer[5][3] , 
        \stage_1_retimer[5][2] , \stage_1_retimer[5][1] , 
        \stage_1_retimer[5][0] }), .in_lower({\stage_1_retimer[7][19] , 
        \stage_1_retimer[7][18] , \stage_1_retimer[7][17] , 
        \stage_1_retimer[7][16] , \stage_1_retimer[7][15] , 
        \stage_1_retimer[7][14] , \stage_1_retimer[7][13] , 
        \stage_1_retimer[7][12] , \stage_1_retimer[7][11] , 
        \stage_1_retimer[7][10] , \stage_1_retimer[7][9] , 
        \stage_1_retimer[7][8] , \stage_1_retimer[7][7] , 
        \stage_1_retimer[7][6] , \stage_1_retimer[7][5] , 
        \stage_1_retimer[7][4] , \stage_1_retimer[7][3] , 
        \stage_1_retimer[7][2] , \stage_1_retimer[7][1] , 
        \stage_1_retimer[7][0] }), .in_control(in_control[8]), .out_upper({
        \stage_2_output[6][19] , \stage_2_output[6][18] , 
        \stage_2_output[6][17] , \stage_2_output[6][16] , 
        \stage_2_output[6][15] , \stage_2_output[6][14] , 
        \stage_2_output[6][13] , \stage_2_output[6][12] , 
        \stage_2_output[6][11] , \stage_2_output[6][10] , 
        \stage_2_output[6][9] , \stage_2_output[6][8] , \stage_2_output[6][7] , 
        \stage_2_output[6][6] , \stage_2_output[6][5] , \stage_2_output[6][4] , 
        \stage_2_output[6][3] , \stage_2_output[6][2] , \stage_2_output[6][1] , 
        \stage_2_output[6][0] }), .out_lower({\stage_2_output[7][19] , 
        \stage_2_output[7][18] , \stage_2_output[7][17] , 
        \stage_2_output[7][16] , \stage_2_output[7][15] , 
        \stage_2_output[7][14] , \stage_2_output[7][13] , 
        \stage_2_output[7][12] , \stage_2_output[7][11] , 
        \stage_2_output[7][10] , \stage_2_output[7][9] , 
        \stage_2_output[7][8] , \stage_2_output[7][7] , \stage_2_output[7][6] , 
        \stage_2_output[7][5] , \stage_2_output[7][4] , \stage_2_output[7][3] , 
        \stage_2_output[7][2] , \stage_2_output[7][1] , \stage_2_output[7][0] }) );
  crossbar_8 u_30_crossbar ( .in_upper({\stage_2_retimer[0][19] , 
        \stage_2_retimer[0][18] , \stage_2_retimer[0][17] , 
        \stage_2_retimer[0][16] , \stage_2_retimer[0][15] , 
        \stage_2_retimer[0][14] , \stage_2_retimer[0][13] , 
        \stage_2_retimer[0][12] , \stage_2_retimer[0][11] , 
        \stage_2_retimer[0][10] , \stage_2_retimer[0][9] , 
        \stage_2_retimer[0][8] , \stage_2_retimer[0][7] , 
        \stage_2_retimer[0][6] , \stage_2_retimer[0][5] , 
        \stage_2_retimer[0][4] , \stage_2_retimer[0][3] , 
        \stage_2_retimer[0][2] , \stage_2_retimer[0][1] , 
        \stage_2_retimer[0][0] }), .in_lower({\stage_2_retimer[2][19] , 
        \stage_2_retimer[2][18] , \stage_2_retimer[2][17] , 
        \stage_2_retimer[2][16] , \stage_2_retimer[2][15] , 
        \stage_2_retimer[2][14] , \stage_2_retimer[2][13] , 
        \stage_2_retimer[2][12] , \stage_2_retimer[2][11] , 
        \stage_2_retimer[2][10] , \stage_2_retimer[2][9] , 
        \stage_2_retimer[2][8] , \stage_2_retimer[2][7] , 
        \stage_2_retimer[2][6] , \stage_2_retimer[2][5] , 
        \stage_2_retimer[2][4] , \stage_2_retimer[2][3] , 
        \stage_2_retimer[2][2] , \stage_2_retimer[2][1] , 
        \stage_2_retimer[2][0] }), .in_control(in_control[7]), .out_upper({
        \stage_3_output[0][19] , \stage_3_output[0][18] , 
        \stage_3_output[0][17] , \stage_3_output[0][16] , 
        \stage_3_output[0][15] , \stage_3_output[0][14] , 
        \stage_3_output[0][13] , \stage_3_output[0][12] , 
        \stage_3_output[0][11] , \stage_3_output[0][10] , 
        \stage_3_output[0][9] , \stage_3_output[0][8] , \stage_3_output[0][7] , 
        \stage_3_output[0][6] , \stage_3_output[0][5] , \stage_3_output[0][4] , 
        \stage_3_output[0][3] , \stage_3_output[0][2] , \stage_3_output[0][1] , 
        \stage_3_output[0][0] }), .out_lower({\stage_3_output[1][19] , 
        \stage_3_output[1][18] , \stage_3_output[1][17] , 
        \stage_3_output[1][16] , \stage_3_output[1][15] , 
        \stage_3_output[1][14] , \stage_3_output[1][13] , 
        \stage_3_output[1][12] , \stage_3_output[1][11] , 
        \stage_3_output[1][10] , \stage_3_output[1][9] , 
        \stage_3_output[1][8] , \stage_3_output[1][7] , \stage_3_output[1][6] , 
        \stage_3_output[1][5] , \stage_3_output[1][4] , \stage_3_output[1][3] , 
        \stage_3_output[1][2] , \stage_3_output[1][1] , \stage_3_output[1][0] }) );
  crossbar_7 u_31_crossbar ( .in_upper({\stage_2_retimer[1][19] , 
        \stage_2_retimer[1][18] , \stage_2_retimer[1][17] , 
        \stage_2_retimer[1][16] , \stage_2_retimer[1][15] , 
        \stage_2_retimer[1][14] , \stage_2_retimer[1][13] , 
        \stage_2_retimer[1][12] , \stage_2_retimer[1][11] , 
        \stage_2_retimer[1][10] , \stage_2_retimer[1][9] , 
        \stage_2_retimer[1][8] , \stage_2_retimer[1][7] , 
        \stage_2_retimer[1][6] , \stage_2_retimer[1][5] , 
        \stage_2_retimer[1][4] , \stage_2_retimer[1][3] , 
        \stage_2_retimer[1][2] , \stage_2_retimer[1][1] , 
        \stage_2_retimer[1][0] }), .in_lower({\stage_2_retimer[3][19] , 
        \stage_2_retimer[3][18] , \stage_2_retimer[3][17] , 
        \stage_2_retimer[3][16] , \stage_2_retimer[3][15] , 
        \stage_2_retimer[3][14] , \stage_2_retimer[3][13] , 
        \stage_2_retimer[3][12] , \stage_2_retimer[3][11] , 
        \stage_2_retimer[3][10] , \stage_2_retimer[3][9] , 
        \stage_2_retimer[3][8] , \stage_2_retimer[3][7] , 
        \stage_2_retimer[3][6] , \stage_2_retimer[3][5] , 
        \stage_2_retimer[3][4] , \stage_2_retimer[3][3] , 
        \stage_2_retimer[3][2] , \stage_2_retimer[3][1] , 
        \stage_2_retimer[3][0] }), .in_control(in_control[6]), .out_upper({
        \stage_3_output[2][19] , \stage_3_output[2][18] , 
        \stage_3_output[2][17] , \stage_3_output[2][16] , 
        \stage_3_output[2][15] , \stage_3_output[2][14] , 
        \stage_3_output[2][13] , \stage_3_output[2][12] , 
        \stage_3_output[2][11] , \stage_3_output[2][10] , 
        \stage_3_output[2][9] , \stage_3_output[2][8] , \stage_3_output[2][7] , 
        \stage_3_output[2][6] , \stage_3_output[2][5] , \stage_3_output[2][4] , 
        \stage_3_output[2][3] , \stage_3_output[2][2] , \stage_3_output[2][1] , 
        \stage_3_output[2][0] }), .out_lower({\stage_3_output[3][19] , 
        \stage_3_output[3][18] , \stage_3_output[3][17] , 
        \stage_3_output[3][16] , \stage_3_output[3][15] , 
        \stage_3_output[3][14] , \stage_3_output[3][13] , 
        \stage_3_output[3][12] , \stage_3_output[3][11] , 
        \stage_3_output[3][10] , \stage_3_output[3][9] , 
        \stage_3_output[3][8] , \stage_3_output[3][7] , \stage_3_output[3][6] , 
        \stage_3_output[3][5] , \stage_3_output[3][4] , \stage_3_output[3][3] , 
        \stage_3_output[3][2] , \stage_3_output[3][1] , \stage_3_output[3][0] }) );
  crossbar_6 u_32_crossbar ( .in_upper({\stage_2_retimer[4][19] , 
        \stage_2_retimer[4][18] , \stage_2_retimer[4][17] , 
        \stage_2_retimer[4][16] , \stage_2_retimer[4][15] , 
        \stage_2_retimer[4][14] , \stage_2_retimer[4][13] , 
        \stage_2_retimer[4][12] , \stage_2_retimer[4][11] , 
        \stage_2_retimer[4][10] , \stage_2_retimer[4][9] , 
        \stage_2_retimer[4][8] , \stage_2_retimer[4][7] , 
        \stage_2_retimer[4][6] , \stage_2_retimer[4][5] , 
        \stage_2_retimer[4][4] , \stage_2_retimer[4][3] , 
        \stage_2_retimer[4][2] , \stage_2_retimer[4][1] , 
        \stage_2_retimer[4][0] }), .in_lower({\stage_2_retimer[6][19] , 
        \stage_2_retimer[6][18] , \stage_2_retimer[6][17] , 
        \stage_2_retimer[6][16] , \stage_2_retimer[6][15] , 
        \stage_2_retimer[6][14] , \stage_2_retimer[6][13] , 
        \stage_2_retimer[6][12] , \stage_2_retimer[6][11] , 
        \stage_2_retimer[6][10] , \stage_2_retimer[6][9] , 
        \stage_2_retimer[6][8] , \stage_2_retimer[6][7] , 
        \stage_2_retimer[6][6] , \stage_2_retimer[6][5] , 
        \stage_2_retimer[6][4] , \stage_2_retimer[6][3] , 
        \stage_2_retimer[6][2] , \stage_2_retimer[6][1] , 
        \stage_2_retimer[6][0] }), .in_control(in_control[5]), .out_upper({
        \stage_3_output[4][19] , \stage_3_output[4][18] , 
        \stage_3_output[4][17] , \stage_3_output[4][16] , 
        \stage_3_output[4][15] , \stage_3_output[4][14] , 
        \stage_3_output[4][13] , \stage_3_output[4][12] , 
        \stage_3_output[4][11] , \stage_3_output[4][10] , 
        \stage_3_output[4][9] , \stage_3_output[4][8] , \stage_3_output[4][7] , 
        \stage_3_output[4][6] , \stage_3_output[4][5] , \stage_3_output[4][4] , 
        \stage_3_output[4][3] , \stage_3_output[4][2] , \stage_3_output[4][1] , 
        \stage_3_output[4][0] }), .out_lower({\stage_3_output[5][19] , 
        \stage_3_output[5][18] , \stage_3_output[5][17] , 
        \stage_3_output[5][16] , \stage_3_output[5][15] , 
        \stage_3_output[5][14] , \stage_3_output[5][13] , 
        \stage_3_output[5][12] , \stage_3_output[5][11] , 
        \stage_3_output[5][10] , \stage_3_output[5][9] , 
        \stage_3_output[5][8] , \stage_3_output[5][7] , \stage_3_output[5][6] , 
        \stage_3_output[5][5] , \stage_3_output[5][4] , \stage_3_output[5][3] , 
        \stage_3_output[5][2] , \stage_3_output[5][1] , \stage_3_output[5][0] }) );
  crossbar_5 u_33_crossbar ( .in_upper({\stage_2_retimer[5][19] , 
        \stage_2_retimer[5][18] , \stage_2_retimer[5][17] , 
        \stage_2_retimer[5][16] , \stage_2_retimer[5][15] , 
        \stage_2_retimer[5][14] , \stage_2_retimer[5][13] , 
        \stage_2_retimer[5][12] , \stage_2_retimer[5][11] , 
        \stage_2_retimer[5][10] , \stage_2_retimer[5][9] , 
        \stage_2_retimer[5][8] , \stage_2_retimer[5][7] , 
        \stage_2_retimer[5][6] , \stage_2_retimer[5][5] , 
        \stage_2_retimer[5][4] , \stage_2_retimer[5][3] , 
        \stage_2_retimer[5][2] , \stage_2_retimer[5][1] , 
        \stage_2_retimer[5][0] }), .in_lower({\stage_2_retimer[7][19] , 
        \stage_2_retimer[7][18] , \stage_2_retimer[7][17] , 
        \stage_2_retimer[7][16] , \stage_2_retimer[7][15] , 
        \stage_2_retimer[7][14] , \stage_2_retimer[7][13] , 
        \stage_2_retimer[7][12] , \stage_2_retimer[7][11] , 
        \stage_2_retimer[7][10] , \stage_2_retimer[7][9] , 
        \stage_2_retimer[7][8] , \stage_2_retimer[7][7] , 
        \stage_2_retimer[7][6] , \stage_2_retimer[7][5] , 
        \stage_2_retimer[7][4] , \stage_2_retimer[7][3] , 
        \stage_2_retimer[7][2] , \stage_2_retimer[7][1] , 
        \stage_2_retimer[7][0] }), .in_control(in_control[4]), .out_upper({
        \stage_3_output[6][19] , \stage_3_output[6][18] , 
        \stage_3_output[6][17] , \stage_3_output[6][16] , 
        \stage_3_output[6][15] , \stage_3_output[6][14] , 
        \stage_3_output[6][13] , \stage_3_output[6][12] , 
        \stage_3_output[6][11] , \stage_3_output[6][10] , 
        \stage_3_output[6][9] , \stage_3_output[6][8] , \stage_3_output[6][7] , 
        \stage_3_output[6][6] , \stage_3_output[6][5] , \stage_3_output[6][4] , 
        \stage_3_output[6][3] , \stage_3_output[6][2] , \stage_3_output[6][1] , 
        \stage_3_output[6][0] }), .out_lower({\stage_3_output[7][19] , 
        \stage_3_output[7][18] , \stage_3_output[7][17] , 
        \stage_3_output[7][16] , \stage_3_output[7][15] , 
        \stage_3_output[7][14] , \stage_3_output[7][13] , 
        \stage_3_output[7][12] , \stage_3_output[7][11] , 
        \stage_3_output[7][10] , \stage_3_output[7][9] , 
        \stage_3_output[7][8] , \stage_3_output[7][7] , \stage_3_output[7][6] , 
        \stage_3_output[7][5] , \stage_3_output[7][4] , \stage_3_output[7][3] , 
        \stage_3_output[7][2] , \stage_3_output[7][1] , \stage_3_output[7][0] }) );
  crossbar_4 u_40_crossbar ( .in_upper({\stage_3_retimer[0][19] , 
        \stage_3_retimer[0][18] , \stage_3_retimer[0][17] , 
        \stage_3_retimer[0][16] , \stage_3_retimer[0][15] , 
        \stage_3_retimer[0][14] , \stage_3_retimer[0][13] , 
        \stage_3_retimer[0][12] , \stage_3_retimer[0][11] , 
        \stage_3_retimer[0][10] , \stage_3_retimer[0][9] , 
        \stage_3_retimer[0][8] , \stage_3_retimer[0][7] , 
        \stage_3_retimer[0][6] , \stage_3_retimer[0][5] , 
        \stage_3_retimer[0][4] , \stage_3_retimer[0][3] , 
        \stage_3_retimer[0][2] , \stage_3_retimer[0][1] , 
        \stage_3_retimer[0][0] }), .in_lower({\stage_3_retimer[4][19] , 
        \stage_3_retimer[4][18] , \stage_3_retimer[4][17] , 
        \stage_3_retimer[4][16] , \stage_3_retimer[4][15] , 
        \stage_3_retimer[4][14] , \stage_3_retimer[4][13] , 
        \stage_3_retimer[4][12] , \stage_3_retimer[4][11] , 
        \stage_3_retimer[4][10] , \stage_3_retimer[4][9] , 
        \stage_3_retimer[4][8] , \stage_3_retimer[4][7] , 
        \stage_3_retimer[4][6] , \stage_3_retimer[4][5] , 
        \stage_3_retimer[4][4] , \stage_3_retimer[4][3] , 
        \stage_3_retimer[4][2] , \stage_3_retimer[4][1] , 
        \stage_3_retimer[4][0] }), .in_control(in_control[3]), .out_upper({
        \stage_4_output[0][19] , \stage_4_output[0][18] , 
        \stage_4_output[0][17] , \stage_4_output[0][16] , 
        \stage_4_output[0][15] , \stage_4_output[0][14] , 
        \stage_4_output[0][13] , \stage_4_output[0][12] , 
        \stage_4_output[0][11] , \stage_4_output[0][10] , 
        \stage_4_output[0][9] , \stage_4_output[0][8] , \stage_4_output[0][7] , 
        \stage_4_output[0][6] , \stage_4_output[0][5] , \stage_4_output[0][4] , 
        \stage_4_output[0][3] , \stage_4_output[0][2] , \stage_4_output[0][1] , 
        \stage_4_output[0][0] }), .out_lower({\stage_4_output[1][19] , 
        \stage_4_output[1][18] , \stage_4_output[1][17] , 
        \stage_4_output[1][16] , \stage_4_output[1][15] , 
        \stage_4_output[1][14] , \stage_4_output[1][13] , 
        \stage_4_output[1][12] , \stage_4_output[1][11] , 
        \stage_4_output[1][10] , \stage_4_output[1][9] , 
        \stage_4_output[1][8] , \stage_4_output[1][7] , \stage_4_output[1][6] , 
        \stage_4_output[1][5] , \stage_4_output[1][4] , \stage_4_output[1][3] , 
        \stage_4_output[1][2] , \stage_4_output[1][1] , \stage_4_output[1][0] }) );
  crossbar_3 u_41_crossbar ( .in_upper({\stage_3_retimer[1][19] , 
        \stage_3_retimer[1][18] , \stage_3_retimer[1][17] , 
        \stage_3_retimer[1][16] , \stage_3_retimer[1][15] , 
        \stage_3_retimer[1][14] , \stage_3_retimer[1][13] , 
        \stage_3_retimer[1][12] , \stage_3_retimer[1][11] , 
        \stage_3_retimer[1][10] , \stage_3_retimer[1][9] , 
        \stage_3_retimer[1][8] , \stage_3_retimer[1][7] , 
        \stage_3_retimer[1][6] , \stage_3_retimer[1][5] , 
        \stage_3_retimer[1][4] , \stage_3_retimer[1][3] , 
        \stage_3_retimer[1][2] , \stage_3_retimer[1][1] , 
        \stage_3_retimer[1][0] }), .in_lower({\stage_3_retimer[5][19] , 
        \stage_3_retimer[5][18] , \stage_3_retimer[5][17] , 
        \stage_3_retimer[5][16] , \stage_3_retimer[5][15] , 
        \stage_3_retimer[5][14] , \stage_3_retimer[5][13] , 
        \stage_3_retimer[5][12] , \stage_3_retimer[5][11] , 
        \stage_3_retimer[5][10] , \stage_3_retimer[5][9] , 
        \stage_3_retimer[5][8] , \stage_3_retimer[5][7] , 
        \stage_3_retimer[5][6] , \stage_3_retimer[5][5] , 
        \stage_3_retimer[5][4] , \stage_3_retimer[5][3] , 
        \stage_3_retimer[5][2] , \stage_3_retimer[5][1] , 
        \stage_3_retimer[5][0] }), .in_control(in_control[2]), .out_upper({
        \stage_4_output[2][19] , \stage_4_output[2][18] , 
        \stage_4_output[2][17] , \stage_4_output[2][16] , 
        \stage_4_output[2][15] , \stage_4_output[2][14] , 
        \stage_4_output[2][13] , \stage_4_output[2][12] , 
        \stage_4_output[2][11] , \stage_4_output[2][10] , 
        \stage_4_output[2][9] , \stage_4_output[2][8] , \stage_4_output[2][7] , 
        \stage_4_output[2][6] , \stage_4_output[2][5] , \stage_4_output[2][4] , 
        \stage_4_output[2][3] , \stage_4_output[2][2] , \stage_4_output[2][1] , 
        \stage_4_output[2][0] }), .out_lower({\stage_4_output[3][19] , 
        \stage_4_output[3][18] , \stage_4_output[3][17] , 
        \stage_4_output[3][16] , \stage_4_output[3][15] , 
        \stage_4_output[3][14] , \stage_4_output[3][13] , 
        \stage_4_output[3][12] , \stage_4_output[3][11] , 
        \stage_4_output[3][10] , \stage_4_output[3][9] , 
        \stage_4_output[3][8] , \stage_4_output[3][7] , \stage_4_output[3][6] , 
        \stage_4_output[3][5] , \stage_4_output[3][4] , \stage_4_output[3][3] , 
        \stage_4_output[3][2] , \stage_4_output[3][1] , \stage_4_output[3][0] }) );
  crossbar_2 u_42_crossbar ( .in_upper({\stage_3_retimer[2][19] , 
        \stage_3_retimer[2][18] , \stage_3_retimer[2][17] , 
        \stage_3_retimer[2][16] , \stage_3_retimer[2][15] , 
        \stage_3_retimer[2][14] , \stage_3_retimer[2][13] , 
        \stage_3_retimer[2][12] , \stage_3_retimer[2][11] , 
        \stage_3_retimer[2][10] , \stage_3_retimer[2][9] , 
        \stage_3_retimer[2][8] , \stage_3_retimer[2][7] , 
        \stage_3_retimer[2][6] , \stage_3_retimer[2][5] , 
        \stage_3_retimer[2][4] , \stage_3_retimer[2][3] , 
        \stage_3_retimer[2][2] , \stage_3_retimer[2][1] , 
        \stage_3_retimer[2][0] }), .in_lower({\stage_3_retimer[6][19] , 
        \stage_3_retimer[6][18] , \stage_3_retimer[6][17] , 
        \stage_3_retimer[6][16] , \stage_3_retimer[6][15] , 
        \stage_3_retimer[6][14] , \stage_3_retimer[6][13] , 
        \stage_3_retimer[6][12] , \stage_3_retimer[6][11] , 
        \stage_3_retimer[6][10] , \stage_3_retimer[6][9] , 
        \stage_3_retimer[6][8] , \stage_3_retimer[6][7] , 
        \stage_3_retimer[6][6] , \stage_3_retimer[6][5] , 
        \stage_3_retimer[6][4] , \stage_3_retimer[6][3] , 
        \stage_3_retimer[6][2] , \stage_3_retimer[6][1] , 
        \stage_3_retimer[6][0] }), .in_control(in_control[1]), .out_upper({
        \stage_4_output[4][19] , \stage_4_output[4][18] , 
        \stage_4_output[4][17] , \stage_4_output[4][16] , 
        \stage_4_output[4][15] , \stage_4_output[4][14] , 
        \stage_4_output[4][13] , \stage_4_output[4][12] , 
        \stage_4_output[4][11] , \stage_4_output[4][10] , 
        \stage_4_output[4][9] , \stage_4_output[4][8] , \stage_4_output[4][7] , 
        \stage_4_output[4][6] , \stage_4_output[4][5] , \stage_4_output[4][4] , 
        \stage_4_output[4][3] , \stage_4_output[4][2] , \stage_4_output[4][1] , 
        \stage_4_output[4][0] }), .out_lower({\stage_4_output[5][19] , 
        \stage_4_output[5][18] , \stage_4_output[5][17] , 
        \stage_4_output[5][16] , \stage_4_output[5][15] , 
        \stage_4_output[5][14] , \stage_4_output[5][13] , 
        \stage_4_output[5][12] , \stage_4_output[5][11] , 
        \stage_4_output[5][10] , \stage_4_output[5][9] , 
        \stage_4_output[5][8] , \stage_4_output[5][7] , \stage_4_output[5][6] , 
        \stage_4_output[5][5] , \stage_4_output[5][4] , \stage_4_output[5][3] , 
        \stage_4_output[5][2] , \stage_4_output[5][1] , \stage_4_output[5][0] }) );
  crossbar_1 u_43_crossbar ( .in_upper({\stage_3_retimer[3][19] , 
        \stage_3_retimer[3][18] , \stage_3_retimer[3][17] , 
        \stage_3_retimer[3][16] , \stage_3_retimer[3][15] , 
        \stage_3_retimer[3][14] , \stage_3_retimer[3][13] , 
        \stage_3_retimer[3][12] , \stage_3_retimer[3][11] , 
        \stage_3_retimer[3][10] , \stage_3_retimer[3][9] , 
        \stage_3_retimer[3][8] , \stage_3_retimer[3][7] , 
        \stage_3_retimer[3][6] , \stage_3_retimer[3][5] , 
        \stage_3_retimer[3][4] , \stage_3_retimer[3][3] , 
        \stage_3_retimer[3][2] , \stage_3_retimer[3][1] , 
        \stage_3_retimer[3][0] }), .in_lower({\stage_3_retimer[7][19] , 
        \stage_3_retimer[7][18] , \stage_3_retimer[7][17] , 
        \stage_3_retimer[7][16] , \stage_3_retimer[7][15] , 
        \stage_3_retimer[7][14] , \stage_3_retimer[7][13] , 
        \stage_3_retimer[7][12] , \stage_3_retimer[7][11] , 
        \stage_3_retimer[7][10] , \stage_3_retimer[7][9] , 
        \stage_3_retimer[7][8] , \stage_3_retimer[7][7] , 
        \stage_3_retimer[7][6] , \stage_3_retimer[7][5] , 
        \stage_3_retimer[7][4] , \stage_3_retimer[7][3] , 
        \stage_3_retimer[7][2] , \stage_3_retimer[7][1] , 
        \stage_3_retimer[7][0] }), .in_control(in_control[0]), .out_upper({
        \stage_4_output[6][19] , \stage_4_output[6][18] , 
        \stage_4_output[6][17] , \stage_4_output[6][16] , 
        \stage_4_output[6][15] , \stage_4_output[6][14] , 
        \stage_4_output[6][13] , \stage_4_output[6][12] , 
        \stage_4_output[6][11] , \stage_4_output[6][10] , 
        \stage_4_output[6][9] , \stage_4_output[6][8] , \stage_4_output[6][7] , 
        \stage_4_output[6][6] , \stage_4_output[6][5] , \stage_4_output[6][4] , 
        \stage_4_output[6][3] , \stage_4_output[6][2] , \stage_4_output[6][1] , 
        \stage_4_output[6][0] }), .out_lower({\stage_4_output[7][19] , 
        \stage_4_output[7][18] , \stage_4_output[7][17] , 
        \stage_4_output[7][16] , \stage_4_output[7][15] , 
        \stage_4_output[7][14] , \stage_4_output[7][13] , 
        \stage_4_output[7][12] , \stage_4_output[7][11] , 
        \stage_4_output[7][10] , \stage_4_output[7][9] , 
        \stage_4_output[7][8] , \stage_4_output[7][7] , \stage_4_output[7][6] , 
        \stage_4_output[7][5] , \stage_4_output[7][4] , \stage_4_output[7][3] , 
        \stage_4_output[7][2] , \stage_4_output[7][1] , \stage_4_output[7][0] }) );
  DFQD1 \stage_0_retimer_reg[7][19]  ( .D(\stage_0_output[7][19] ), .CP(clk), 
        .Q(\stage_0_retimer[7][19] ) );
  DFQD1 \stage_0_retimer_reg[7][18]  ( .D(\stage_0_output[7][18] ), .CP(clk), 
        .Q(\stage_0_retimer[7][18] ) );
  DFQD1 \stage_0_retimer_reg[7][17]  ( .D(\stage_0_output[7][17] ), .CP(clk), 
        .Q(\stage_0_retimer[7][17] ) );
  DFQD1 \stage_0_retimer_reg[7][16]  ( .D(\stage_0_output[7][16] ), .CP(clk), 
        .Q(\stage_0_retimer[7][16] ) );
  DFQD1 \stage_0_retimer_reg[7][15]  ( .D(\stage_0_output[7][15] ), .CP(clk), 
        .Q(\stage_0_retimer[7][15] ) );
  DFQD1 \stage_0_retimer_reg[7][14]  ( .D(\stage_0_output[7][14] ), .CP(clk), 
        .Q(\stage_0_retimer[7][14] ) );
  DFQD1 \stage_0_retimer_reg[7][13]  ( .D(\stage_0_output[7][13] ), .CP(clk), 
        .Q(\stage_0_retimer[7][13] ) );
  DFQD1 \stage_0_retimer_reg[7][12]  ( .D(\stage_0_output[7][12] ), .CP(clk), 
        .Q(\stage_0_retimer[7][12] ) );
  DFQD1 \stage_0_retimer_reg[7][11]  ( .D(\stage_0_output[7][11] ), .CP(clk), 
        .Q(\stage_0_retimer[7][11] ) );
  DFQD1 \stage_0_retimer_reg[7][10]  ( .D(\stage_0_output[7][10] ), .CP(clk), 
        .Q(\stage_0_retimer[7][10] ) );
  DFQD1 \stage_0_retimer_reg[7][9]  ( .D(\stage_0_output[7][9] ), .CP(clk), 
        .Q(\stage_0_retimer[7][9] ) );
  DFQD1 \stage_0_retimer_reg[7][8]  ( .D(\stage_0_output[7][8] ), .CP(clk), 
        .Q(\stage_0_retimer[7][8] ) );
  DFQD1 \stage_0_retimer_reg[7][7]  ( .D(\stage_0_output[7][7] ), .CP(clk), 
        .Q(\stage_0_retimer[7][7] ) );
  DFQD1 \stage_0_retimer_reg[7][6]  ( .D(\stage_0_output[7][6] ), .CP(clk), 
        .Q(\stage_0_retimer[7][6] ) );
  DFQD1 \stage_0_retimer_reg[7][5]  ( .D(\stage_0_output[7][5] ), .CP(clk), 
        .Q(\stage_0_retimer[7][5] ) );
  DFQD1 \stage_0_retimer_reg[7][4]  ( .D(\stage_0_output[7][4] ), .CP(clk), 
        .Q(\stage_0_retimer[7][4] ) );
  DFQD1 \stage_0_retimer_reg[7][3]  ( .D(\stage_0_output[7][3] ), .CP(clk), 
        .Q(\stage_0_retimer[7][3] ) );
  DFQD1 \stage_0_retimer_reg[7][2]  ( .D(\stage_0_output[7][2] ), .CP(clk), 
        .Q(\stage_0_retimer[7][2] ) );
  DFQD1 \stage_0_retimer_reg[7][1]  ( .D(\stage_0_output[7][1] ), .CP(clk), 
        .Q(\stage_0_retimer[7][1] ) );
  DFQD1 \stage_0_retimer_reg[7][0]  ( .D(\stage_0_output[7][0] ), .CP(clk), 
        .Q(\stage_0_retimer[7][0] ) );
  DFQD1 \stage_0_retimer_reg[6][19]  ( .D(\stage_0_output[6][19] ), .CP(clk), 
        .Q(\stage_0_retimer[6][19] ) );
  DFQD1 \stage_0_retimer_reg[6][18]  ( .D(\stage_0_output[6][18] ), .CP(clk), 
        .Q(\stage_0_retimer[6][18] ) );
  DFQD1 \stage_0_retimer_reg[6][17]  ( .D(\stage_0_output[6][17] ), .CP(clk), 
        .Q(\stage_0_retimer[6][17] ) );
  DFQD1 \stage_0_retimer_reg[6][16]  ( .D(\stage_0_output[6][16] ), .CP(clk), 
        .Q(\stage_0_retimer[6][16] ) );
  DFQD1 \stage_0_retimer_reg[6][15]  ( .D(\stage_0_output[6][15] ), .CP(clk), 
        .Q(\stage_0_retimer[6][15] ) );
  DFQD1 \stage_0_retimer_reg[6][14]  ( .D(\stage_0_output[6][14] ), .CP(clk), 
        .Q(\stage_0_retimer[6][14] ) );
  DFQD1 \stage_0_retimer_reg[6][13]  ( .D(\stage_0_output[6][13] ), .CP(clk), 
        .Q(\stage_0_retimer[6][13] ) );
  DFQD1 \stage_0_retimer_reg[6][12]  ( .D(\stage_0_output[6][12] ), .CP(clk), 
        .Q(\stage_0_retimer[6][12] ) );
  DFQD1 \stage_0_retimer_reg[6][11]  ( .D(\stage_0_output[6][11] ), .CP(clk), 
        .Q(\stage_0_retimer[6][11] ) );
  DFQD1 \stage_0_retimer_reg[6][10]  ( .D(\stage_0_output[6][10] ), .CP(clk), 
        .Q(\stage_0_retimer[6][10] ) );
  DFQD1 \stage_0_retimer_reg[6][9]  ( .D(\stage_0_output[6][9] ), .CP(clk), 
        .Q(\stage_0_retimer[6][9] ) );
  DFQD1 \stage_0_retimer_reg[6][8]  ( .D(\stage_0_output[6][8] ), .CP(clk), 
        .Q(\stage_0_retimer[6][8] ) );
  DFQD1 \stage_0_retimer_reg[6][7]  ( .D(\stage_0_output[6][7] ), .CP(clk), 
        .Q(\stage_0_retimer[6][7] ) );
  DFQD1 \stage_0_retimer_reg[6][6]  ( .D(\stage_0_output[6][6] ), .CP(clk), 
        .Q(\stage_0_retimer[6][6] ) );
  DFQD1 \stage_0_retimer_reg[6][5]  ( .D(\stage_0_output[6][5] ), .CP(clk), 
        .Q(\stage_0_retimer[6][5] ) );
  DFQD1 \stage_0_retimer_reg[6][4]  ( .D(\stage_0_output[6][4] ), .CP(clk), 
        .Q(\stage_0_retimer[6][4] ) );
  DFQD1 \stage_0_retimer_reg[6][3]  ( .D(\stage_0_output[6][3] ), .CP(clk), 
        .Q(\stage_0_retimer[6][3] ) );
  DFQD1 \stage_0_retimer_reg[6][2]  ( .D(\stage_0_output[6][2] ), .CP(clk), 
        .Q(\stage_0_retimer[6][2] ) );
  DFQD1 \stage_0_retimer_reg[6][1]  ( .D(\stage_0_output[6][1] ), .CP(clk), 
        .Q(\stage_0_retimer[6][1] ) );
  DFQD1 \stage_0_retimer_reg[6][0]  ( .D(\stage_0_output[6][0] ), .CP(clk), 
        .Q(\stage_0_retimer[6][0] ) );
  DFQD1 \stage_0_retimer_reg[5][19]  ( .D(\stage_0_output[5][19] ), .CP(clk), 
        .Q(\stage_0_retimer[5][19] ) );
  DFQD1 \stage_0_retimer_reg[5][18]  ( .D(\stage_0_output[5][18] ), .CP(clk), 
        .Q(\stage_0_retimer[5][18] ) );
  DFQD1 \stage_0_retimer_reg[5][17]  ( .D(\stage_0_output[5][17] ), .CP(clk), 
        .Q(\stage_0_retimer[5][17] ) );
  DFQD1 \stage_0_retimer_reg[5][16]  ( .D(\stage_0_output[5][16] ), .CP(clk), 
        .Q(\stage_0_retimer[5][16] ) );
  DFQD1 \stage_0_retimer_reg[5][15]  ( .D(\stage_0_output[5][15] ), .CP(clk), 
        .Q(\stage_0_retimer[5][15] ) );
  DFQD1 \stage_0_retimer_reg[5][14]  ( .D(\stage_0_output[5][14] ), .CP(clk), 
        .Q(\stage_0_retimer[5][14] ) );
  DFQD1 \stage_0_retimer_reg[5][13]  ( .D(\stage_0_output[5][13] ), .CP(clk), 
        .Q(\stage_0_retimer[5][13] ) );
  DFQD1 \stage_0_retimer_reg[5][12]  ( .D(\stage_0_output[5][12] ), .CP(clk), 
        .Q(\stage_0_retimer[5][12] ) );
  DFQD1 \stage_0_retimer_reg[5][11]  ( .D(\stage_0_output[5][11] ), .CP(clk), 
        .Q(\stage_0_retimer[5][11] ) );
  DFQD1 \stage_0_retimer_reg[5][10]  ( .D(\stage_0_output[5][10] ), .CP(clk), 
        .Q(\stage_0_retimer[5][10] ) );
  DFQD1 \stage_0_retimer_reg[5][9]  ( .D(\stage_0_output[5][9] ), .CP(clk), 
        .Q(\stage_0_retimer[5][9] ) );
  DFQD1 \stage_0_retimer_reg[5][8]  ( .D(\stage_0_output[5][8] ), .CP(clk), 
        .Q(\stage_0_retimer[5][8] ) );
  DFQD1 \stage_0_retimer_reg[5][7]  ( .D(\stage_0_output[5][7] ), .CP(clk), 
        .Q(\stage_0_retimer[5][7] ) );
  DFQD1 \stage_0_retimer_reg[5][6]  ( .D(\stage_0_output[5][6] ), .CP(clk), 
        .Q(\stage_0_retimer[5][6] ) );
  DFQD1 \stage_0_retimer_reg[5][5]  ( .D(\stage_0_output[5][5] ), .CP(clk), 
        .Q(\stage_0_retimer[5][5] ) );
  DFQD1 \stage_0_retimer_reg[5][4]  ( .D(\stage_0_output[5][4] ), .CP(clk), 
        .Q(\stage_0_retimer[5][4] ) );
  DFQD1 \stage_0_retimer_reg[5][3]  ( .D(\stage_0_output[5][3] ), .CP(clk), 
        .Q(\stage_0_retimer[5][3] ) );
  DFQD1 \stage_0_retimer_reg[5][2]  ( .D(\stage_0_output[5][2] ), .CP(clk), 
        .Q(\stage_0_retimer[5][2] ) );
  DFQD1 \stage_0_retimer_reg[5][1]  ( .D(\stage_0_output[5][1] ), .CP(clk), 
        .Q(\stage_0_retimer[5][1] ) );
  DFQD1 \stage_0_retimer_reg[5][0]  ( .D(\stage_0_output[5][0] ), .CP(clk), 
        .Q(\stage_0_retimer[5][0] ) );
  DFQD1 \stage_0_retimer_reg[4][19]  ( .D(\stage_0_output[4][19] ), .CP(clk), 
        .Q(\stage_0_retimer[4][19] ) );
  DFQD1 \stage_0_retimer_reg[4][18]  ( .D(\stage_0_output[4][18] ), .CP(clk), 
        .Q(\stage_0_retimer[4][18] ) );
  DFQD1 \stage_0_retimer_reg[4][17]  ( .D(\stage_0_output[4][17] ), .CP(clk), 
        .Q(\stage_0_retimer[4][17] ) );
  DFQD1 \stage_0_retimer_reg[4][16]  ( .D(\stage_0_output[4][16] ), .CP(clk), 
        .Q(\stage_0_retimer[4][16] ) );
  DFQD1 \stage_0_retimer_reg[4][15]  ( .D(\stage_0_output[4][15] ), .CP(clk), 
        .Q(\stage_0_retimer[4][15] ) );
  DFQD1 \stage_0_retimer_reg[4][14]  ( .D(\stage_0_output[4][14] ), .CP(clk), 
        .Q(\stage_0_retimer[4][14] ) );
  DFQD1 \stage_0_retimer_reg[4][13]  ( .D(\stage_0_output[4][13] ), .CP(clk), 
        .Q(\stage_0_retimer[4][13] ) );
  DFQD1 \stage_0_retimer_reg[4][12]  ( .D(\stage_0_output[4][12] ), .CP(clk), 
        .Q(\stage_0_retimer[4][12] ) );
  DFQD1 \stage_0_retimer_reg[4][11]  ( .D(\stage_0_output[4][11] ), .CP(clk), 
        .Q(\stage_0_retimer[4][11] ) );
  DFQD1 \stage_0_retimer_reg[4][10]  ( .D(\stage_0_output[4][10] ), .CP(clk), 
        .Q(\stage_0_retimer[4][10] ) );
  DFQD1 \stage_0_retimer_reg[4][9]  ( .D(\stage_0_output[4][9] ), .CP(clk), 
        .Q(\stage_0_retimer[4][9] ) );
  DFQD1 \stage_0_retimer_reg[4][8]  ( .D(\stage_0_output[4][8] ), .CP(clk), 
        .Q(\stage_0_retimer[4][8] ) );
  DFQD1 \stage_0_retimer_reg[4][7]  ( .D(\stage_0_output[4][7] ), .CP(clk), 
        .Q(\stage_0_retimer[4][7] ) );
  DFQD1 \stage_0_retimer_reg[4][6]  ( .D(\stage_0_output[4][6] ), .CP(clk), 
        .Q(\stage_0_retimer[4][6] ) );
  DFQD1 \stage_0_retimer_reg[4][5]  ( .D(\stage_0_output[4][5] ), .CP(clk), 
        .Q(\stage_0_retimer[4][5] ) );
  DFQD1 \stage_0_retimer_reg[4][4]  ( .D(\stage_0_output[4][4] ), .CP(clk), 
        .Q(\stage_0_retimer[4][4] ) );
  DFQD1 \stage_0_retimer_reg[4][3]  ( .D(\stage_0_output[4][3] ), .CP(clk), 
        .Q(\stage_0_retimer[4][3] ) );
  DFQD1 \stage_0_retimer_reg[4][2]  ( .D(\stage_0_output[4][2] ), .CP(clk), 
        .Q(\stage_0_retimer[4][2] ) );
  DFQD1 \stage_0_retimer_reg[4][1]  ( .D(\stage_0_output[4][1] ), .CP(clk), 
        .Q(\stage_0_retimer[4][1] ) );
  DFQD1 \stage_0_retimer_reg[4][0]  ( .D(\stage_0_output[4][0] ), .CP(clk), 
        .Q(\stage_0_retimer[4][0] ) );
  DFQD1 \stage_0_retimer_reg[3][19]  ( .D(\stage_0_output[3][19] ), .CP(clk), 
        .Q(\stage_0_retimer[3][19] ) );
  DFQD1 \stage_0_retimer_reg[3][18]  ( .D(\stage_0_output[3][18] ), .CP(clk), 
        .Q(\stage_0_retimer[3][18] ) );
  DFQD1 \stage_0_retimer_reg[3][17]  ( .D(\stage_0_output[3][17] ), .CP(clk), 
        .Q(\stage_0_retimer[3][17] ) );
  DFQD1 \stage_0_retimer_reg[3][16]  ( .D(\stage_0_output[3][16] ), .CP(clk), 
        .Q(\stage_0_retimer[3][16] ) );
  DFQD1 \stage_0_retimer_reg[3][15]  ( .D(\stage_0_output[3][15] ), .CP(clk), 
        .Q(\stage_0_retimer[3][15] ) );
  DFQD1 \stage_0_retimer_reg[3][14]  ( .D(\stage_0_output[3][14] ), .CP(clk), 
        .Q(\stage_0_retimer[3][14] ) );
  DFQD1 \stage_0_retimer_reg[3][13]  ( .D(\stage_0_output[3][13] ), .CP(clk), 
        .Q(\stage_0_retimer[3][13] ) );
  DFQD1 \stage_0_retimer_reg[3][12]  ( .D(\stage_0_output[3][12] ), .CP(clk), 
        .Q(\stage_0_retimer[3][12] ) );
  DFQD1 \stage_0_retimer_reg[3][11]  ( .D(\stage_0_output[3][11] ), .CP(clk), 
        .Q(\stage_0_retimer[3][11] ) );
  DFQD1 \stage_0_retimer_reg[3][10]  ( .D(\stage_0_output[3][10] ), .CP(clk), 
        .Q(\stage_0_retimer[3][10] ) );
  DFQD1 \stage_0_retimer_reg[3][9]  ( .D(\stage_0_output[3][9] ), .CP(clk), 
        .Q(\stage_0_retimer[3][9] ) );
  DFQD1 \stage_0_retimer_reg[3][8]  ( .D(\stage_0_output[3][8] ), .CP(clk), 
        .Q(\stage_0_retimer[3][8] ) );
  DFQD1 \stage_0_retimer_reg[3][7]  ( .D(\stage_0_output[3][7] ), .CP(clk), 
        .Q(\stage_0_retimer[3][7] ) );
  DFQD1 \stage_0_retimer_reg[3][6]  ( .D(\stage_0_output[3][6] ), .CP(clk), 
        .Q(\stage_0_retimer[3][6] ) );
  DFQD1 \stage_0_retimer_reg[3][5]  ( .D(\stage_0_output[3][5] ), .CP(clk), 
        .Q(\stage_0_retimer[3][5] ) );
  DFQD1 \stage_0_retimer_reg[3][4]  ( .D(\stage_0_output[3][4] ), .CP(clk), 
        .Q(\stage_0_retimer[3][4] ) );
  DFQD1 \stage_0_retimer_reg[3][3]  ( .D(\stage_0_output[3][3] ), .CP(clk), 
        .Q(\stage_0_retimer[3][3] ) );
  DFQD1 \stage_0_retimer_reg[3][2]  ( .D(\stage_0_output[3][2] ), .CP(clk), 
        .Q(\stage_0_retimer[3][2] ) );
  DFQD1 \stage_0_retimer_reg[3][1]  ( .D(\stage_0_output[3][1] ), .CP(clk), 
        .Q(\stage_0_retimer[3][1] ) );
  DFQD1 \stage_0_retimer_reg[3][0]  ( .D(\stage_0_output[3][0] ), .CP(clk), 
        .Q(\stage_0_retimer[3][0] ) );
  DFQD1 \stage_0_retimer_reg[2][19]  ( .D(\stage_0_output[2][19] ), .CP(clk), 
        .Q(\stage_0_retimer[2][19] ) );
  DFQD1 \stage_0_retimer_reg[2][18]  ( .D(\stage_0_output[2][18] ), .CP(clk), 
        .Q(\stage_0_retimer[2][18] ) );
  DFQD1 \stage_0_retimer_reg[2][17]  ( .D(\stage_0_output[2][17] ), .CP(clk), 
        .Q(\stage_0_retimer[2][17] ) );
  DFQD1 \stage_0_retimer_reg[2][16]  ( .D(\stage_0_output[2][16] ), .CP(clk), 
        .Q(\stage_0_retimer[2][16] ) );
  DFQD1 \stage_0_retimer_reg[2][15]  ( .D(\stage_0_output[2][15] ), .CP(clk), 
        .Q(\stage_0_retimer[2][15] ) );
  DFQD1 \stage_0_retimer_reg[2][14]  ( .D(\stage_0_output[2][14] ), .CP(clk), 
        .Q(\stage_0_retimer[2][14] ) );
  DFQD1 \stage_0_retimer_reg[2][13]  ( .D(\stage_0_output[2][13] ), .CP(clk), 
        .Q(\stage_0_retimer[2][13] ) );
  DFQD1 \stage_0_retimer_reg[2][12]  ( .D(\stage_0_output[2][12] ), .CP(clk), 
        .Q(\stage_0_retimer[2][12] ) );
  DFQD1 \stage_0_retimer_reg[2][11]  ( .D(\stage_0_output[2][11] ), .CP(clk), 
        .Q(\stage_0_retimer[2][11] ) );
  DFQD1 \stage_0_retimer_reg[2][10]  ( .D(\stage_0_output[2][10] ), .CP(clk), 
        .Q(\stage_0_retimer[2][10] ) );
  DFQD1 \stage_0_retimer_reg[2][9]  ( .D(\stage_0_output[2][9] ), .CP(clk), 
        .Q(\stage_0_retimer[2][9] ) );
  DFQD1 \stage_0_retimer_reg[2][8]  ( .D(\stage_0_output[2][8] ), .CP(clk), 
        .Q(\stage_0_retimer[2][8] ) );
  DFQD1 \stage_0_retimer_reg[2][7]  ( .D(\stage_0_output[2][7] ), .CP(clk), 
        .Q(\stage_0_retimer[2][7] ) );
  DFQD1 \stage_0_retimer_reg[2][6]  ( .D(\stage_0_output[2][6] ), .CP(clk), 
        .Q(\stage_0_retimer[2][6] ) );
  DFQD1 \stage_0_retimer_reg[2][5]  ( .D(\stage_0_output[2][5] ), .CP(clk), 
        .Q(\stage_0_retimer[2][5] ) );
  DFQD1 \stage_0_retimer_reg[2][4]  ( .D(\stage_0_output[2][4] ), .CP(clk), 
        .Q(\stage_0_retimer[2][4] ) );
  DFQD1 \stage_0_retimer_reg[2][3]  ( .D(\stage_0_output[2][3] ), .CP(clk), 
        .Q(\stage_0_retimer[2][3] ) );
  DFQD1 \stage_0_retimer_reg[2][2]  ( .D(\stage_0_output[2][2] ), .CP(clk), 
        .Q(\stage_0_retimer[2][2] ) );
  DFQD1 \stage_0_retimer_reg[2][1]  ( .D(\stage_0_output[2][1] ), .CP(clk), 
        .Q(\stage_0_retimer[2][1] ) );
  DFQD1 \stage_0_retimer_reg[2][0]  ( .D(\stage_0_output[2][0] ), .CP(clk), 
        .Q(\stage_0_retimer[2][0] ) );
  DFQD1 \stage_0_retimer_reg[1][19]  ( .D(\stage_0_output[1][19] ), .CP(clk), 
        .Q(\stage_0_retimer[1][19] ) );
  DFQD1 \stage_0_retimer_reg[1][18]  ( .D(\stage_0_output[1][18] ), .CP(clk), 
        .Q(\stage_0_retimer[1][18] ) );
  DFQD1 \stage_0_retimer_reg[1][17]  ( .D(\stage_0_output[1][17] ), .CP(clk), 
        .Q(\stage_0_retimer[1][17] ) );
  DFQD1 \stage_0_retimer_reg[1][16]  ( .D(\stage_0_output[1][16] ), .CP(clk), 
        .Q(\stage_0_retimer[1][16] ) );
  DFQD1 \stage_0_retimer_reg[1][15]  ( .D(\stage_0_output[1][15] ), .CP(clk), 
        .Q(\stage_0_retimer[1][15] ) );
  DFQD1 \stage_0_retimer_reg[1][14]  ( .D(\stage_0_output[1][14] ), .CP(clk), 
        .Q(\stage_0_retimer[1][14] ) );
  DFQD1 \stage_0_retimer_reg[1][13]  ( .D(\stage_0_output[1][13] ), .CP(clk), 
        .Q(\stage_0_retimer[1][13] ) );
  DFQD1 \stage_0_retimer_reg[1][12]  ( .D(\stage_0_output[1][12] ), .CP(clk), 
        .Q(\stage_0_retimer[1][12] ) );
  DFQD1 \stage_0_retimer_reg[1][11]  ( .D(\stage_0_output[1][11] ), .CP(clk), 
        .Q(\stage_0_retimer[1][11] ) );
  DFQD1 \stage_0_retimer_reg[1][10]  ( .D(\stage_0_output[1][10] ), .CP(clk), 
        .Q(\stage_0_retimer[1][10] ) );
  DFQD1 \stage_0_retimer_reg[1][9]  ( .D(\stage_0_output[1][9] ), .CP(clk), 
        .Q(\stage_0_retimer[1][9] ) );
  DFQD1 \stage_0_retimer_reg[1][8]  ( .D(\stage_0_output[1][8] ), .CP(clk), 
        .Q(\stage_0_retimer[1][8] ) );
  DFQD1 \stage_0_retimer_reg[1][7]  ( .D(\stage_0_output[1][7] ), .CP(clk), 
        .Q(\stage_0_retimer[1][7] ) );
  DFQD1 \stage_0_retimer_reg[1][6]  ( .D(\stage_0_output[1][6] ), .CP(clk), 
        .Q(\stage_0_retimer[1][6] ) );
  DFQD1 \stage_0_retimer_reg[1][5]  ( .D(\stage_0_output[1][5] ), .CP(clk), 
        .Q(\stage_0_retimer[1][5] ) );
  DFQD1 \stage_0_retimer_reg[1][4]  ( .D(\stage_0_output[1][4] ), .CP(clk), 
        .Q(\stage_0_retimer[1][4] ) );
  DFQD1 \stage_0_retimer_reg[1][3]  ( .D(\stage_0_output[1][3] ), .CP(clk), 
        .Q(\stage_0_retimer[1][3] ) );
  DFQD1 \stage_0_retimer_reg[1][2]  ( .D(\stage_0_output[1][2] ), .CP(clk), 
        .Q(\stage_0_retimer[1][2] ) );
  DFQD1 \stage_0_retimer_reg[1][1]  ( .D(\stage_0_output[1][1] ), .CP(clk), 
        .Q(\stage_0_retimer[1][1] ) );
  DFQD1 \stage_0_retimer_reg[1][0]  ( .D(\stage_0_output[1][0] ), .CP(clk), 
        .Q(\stage_0_retimer[1][0] ) );
  DFQD1 \stage_0_retimer_reg[0][19]  ( .D(\stage_0_output[0][19] ), .CP(clk), 
        .Q(\stage_0_retimer[0][19] ) );
  DFQD1 \stage_0_retimer_reg[0][18]  ( .D(\stage_0_output[0][18] ), .CP(clk), 
        .Q(\stage_0_retimer[0][18] ) );
  DFQD1 \stage_0_retimer_reg[0][17]  ( .D(\stage_0_output[0][17] ), .CP(clk), 
        .Q(\stage_0_retimer[0][17] ) );
  DFQD1 \stage_0_retimer_reg[0][16]  ( .D(\stage_0_output[0][16] ), .CP(clk), 
        .Q(\stage_0_retimer[0][16] ) );
  DFQD1 \stage_0_retimer_reg[0][15]  ( .D(\stage_0_output[0][15] ), .CP(clk), 
        .Q(\stage_0_retimer[0][15] ) );
  DFQD1 \stage_0_retimer_reg[0][14]  ( .D(\stage_0_output[0][14] ), .CP(clk), 
        .Q(\stage_0_retimer[0][14] ) );
  DFQD1 \stage_0_retimer_reg[0][13]  ( .D(\stage_0_output[0][13] ), .CP(clk), 
        .Q(\stage_0_retimer[0][13] ) );
  DFQD1 \stage_0_retimer_reg[0][12]  ( .D(\stage_0_output[0][12] ), .CP(clk), 
        .Q(\stage_0_retimer[0][12] ) );
  DFQD1 \stage_0_retimer_reg[0][11]  ( .D(\stage_0_output[0][11] ), .CP(clk), 
        .Q(\stage_0_retimer[0][11] ) );
  DFQD1 \stage_0_retimer_reg[0][10]  ( .D(\stage_0_output[0][10] ), .CP(clk), 
        .Q(\stage_0_retimer[0][10] ) );
  DFQD1 \stage_0_retimer_reg[0][9]  ( .D(\stage_0_output[0][9] ), .CP(clk), 
        .Q(\stage_0_retimer[0][9] ) );
  DFQD1 \stage_0_retimer_reg[0][8]  ( .D(\stage_0_output[0][8] ), .CP(clk), 
        .Q(\stage_0_retimer[0][8] ) );
  DFQD1 \stage_0_retimer_reg[0][7]  ( .D(\stage_0_output[0][7] ), .CP(clk), 
        .Q(\stage_0_retimer[0][7] ) );
  DFQD1 \stage_0_retimer_reg[0][6]  ( .D(\stage_0_output[0][6] ), .CP(clk), 
        .Q(\stage_0_retimer[0][6] ) );
  DFQD1 \stage_0_retimer_reg[0][5]  ( .D(\stage_0_output[0][5] ), .CP(clk), 
        .Q(\stage_0_retimer[0][5] ) );
  DFQD1 \stage_0_retimer_reg[0][4]  ( .D(\stage_0_output[0][4] ), .CP(clk), 
        .Q(\stage_0_retimer[0][4] ) );
  DFQD1 \stage_0_retimer_reg[0][3]  ( .D(\stage_0_output[0][3] ), .CP(clk), 
        .Q(\stage_0_retimer[0][3] ) );
  DFQD1 \stage_0_retimer_reg[0][2]  ( .D(\stage_0_output[0][2] ), .CP(clk), 
        .Q(\stage_0_retimer[0][2] ) );
  DFQD1 \stage_0_retimer_reg[0][1]  ( .D(\stage_0_output[0][1] ), .CP(clk), 
        .Q(\stage_0_retimer[0][1] ) );
  DFQD1 \stage_0_retimer_reg[0][0]  ( .D(\stage_0_output[0][0] ), .CP(clk), 
        .Q(\stage_0_retimer[0][0] ) );
  DFQD1 \stage_1_retimer_reg[7][19]  ( .D(\stage_1_output[7][19] ), .CP(clk), 
        .Q(\stage_1_retimer[7][19] ) );
  DFQD1 \stage_1_retimer_reg[7][18]  ( .D(\stage_1_output[7][18] ), .CP(clk), 
        .Q(\stage_1_retimer[7][18] ) );
  DFQD1 \stage_1_retimer_reg[7][17]  ( .D(\stage_1_output[7][17] ), .CP(clk), 
        .Q(\stage_1_retimer[7][17] ) );
  DFQD1 \stage_1_retimer_reg[7][16]  ( .D(\stage_1_output[7][16] ), .CP(clk), 
        .Q(\stage_1_retimer[7][16] ) );
  DFQD1 \stage_1_retimer_reg[7][15]  ( .D(\stage_1_output[7][15] ), .CP(clk), 
        .Q(\stage_1_retimer[7][15] ) );
  DFQD1 \stage_1_retimer_reg[7][14]  ( .D(\stage_1_output[7][14] ), .CP(clk), 
        .Q(\stage_1_retimer[7][14] ) );
  DFQD1 \stage_1_retimer_reg[7][13]  ( .D(\stage_1_output[7][13] ), .CP(clk), 
        .Q(\stage_1_retimer[7][13] ) );
  DFQD1 \stage_1_retimer_reg[7][12]  ( .D(\stage_1_output[7][12] ), .CP(clk), 
        .Q(\stage_1_retimer[7][12] ) );
  DFQD1 \stage_1_retimer_reg[7][11]  ( .D(\stage_1_output[7][11] ), .CP(clk), 
        .Q(\stage_1_retimer[7][11] ) );
  DFQD1 \stage_1_retimer_reg[7][10]  ( .D(\stage_1_output[7][10] ), .CP(clk), 
        .Q(\stage_1_retimer[7][10] ) );
  DFQD1 \stage_1_retimer_reg[7][9]  ( .D(\stage_1_output[7][9] ), .CP(clk), 
        .Q(\stage_1_retimer[7][9] ) );
  DFQD1 \stage_1_retimer_reg[7][8]  ( .D(\stage_1_output[7][8] ), .CP(clk), 
        .Q(\stage_1_retimer[7][8] ) );
  DFQD1 \stage_1_retimer_reg[7][7]  ( .D(\stage_1_output[7][7] ), .CP(clk), 
        .Q(\stage_1_retimer[7][7] ) );
  DFQD1 \stage_1_retimer_reg[7][6]  ( .D(\stage_1_output[7][6] ), .CP(clk), 
        .Q(\stage_1_retimer[7][6] ) );
  DFQD1 \stage_1_retimer_reg[7][5]  ( .D(\stage_1_output[7][5] ), .CP(clk), 
        .Q(\stage_1_retimer[7][5] ) );
  DFQD1 \stage_1_retimer_reg[7][4]  ( .D(\stage_1_output[7][4] ), .CP(clk), 
        .Q(\stage_1_retimer[7][4] ) );
  DFQD1 \stage_1_retimer_reg[7][3]  ( .D(\stage_1_output[7][3] ), .CP(clk), 
        .Q(\stage_1_retimer[7][3] ) );
  DFQD1 \stage_1_retimer_reg[7][2]  ( .D(\stage_1_output[7][2] ), .CP(clk), 
        .Q(\stage_1_retimer[7][2] ) );
  DFQD1 \stage_1_retimer_reg[7][1]  ( .D(\stage_1_output[7][1] ), .CP(clk), 
        .Q(\stage_1_retimer[7][1] ) );
  DFQD1 \stage_1_retimer_reg[7][0]  ( .D(\stage_1_output[7][0] ), .CP(clk), 
        .Q(\stage_1_retimer[7][0] ) );
  DFQD1 \stage_1_retimer_reg[6][19]  ( .D(\stage_1_output[6][19] ), .CP(clk), 
        .Q(\stage_1_retimer[6][19] ) );
  DFQD1 \stage_1_retimer_reg[6][18]  ( .D(\stage_1_output[6][18] ), .CP(clk), 
        .Q(\stage_1_retimer[6][18] ) );
  DFQD1 \stage_1_retimer_reg[6][17]  ( .D(\stage_1_output[6][17] ), .CP(clk), 
        .Q(\stage_1_retimer[6][17] ) );
  DFQD1 \stage_1_retimer_reg[6][16]  ( .D(\stage_1_output[6][16] ), .CP(clk), 
        .Q(\stage_1_retimer[6][16] ) );
  DFQD1 \stage_1_retimer_reg[6][15]  ( .D(\stage_1_output[6][15] ), .CP(clk), 
        .Q(\stage_1_retimer[6][15] ) );
  DFQD1 \stage_1_retimer_reg[6][14]  ( .D(\stage_1_output[6][14] ), .CP(clk), 
        .Q(\stage_1_retimer[6][14] ) );
  DFQD1 \stage_1_retimer_reg[6][13]  ( .D(\stage_1_output[6][13] ), .CP(clk), 
        .Q(\stage_1_retimer[6][13] ) );
  DFQD1 \stage_1_retimer_reg[6][12]  ( .D(\stage_1_output[6][12] ), .CP(clk), 
        .Q(\stage_1_retimer[6][12] ) );
  DFQD1 \stage_1_retimer_reg[6][11]  ( .D(\stage_1_output[6][11] ), .CP(clk), 
        .Q(\stage_1_retimer[6][11] ) );
  DFQD1 \stage_1_retimer_reg[6][10]  ( .D(\stage_1_output[6][10] ), .CP(clk), 
        .Q(\stage_1_retimer[6][10] ) );
  DFQD1 \stage_1_retimer_reg[6][9]  ( .D(\stage_1_output[6][9] ), .CP(clk), 
        .Q(\stage_1_retimer[6][9] ) );
  DFQD1 \stage_1_retimer_reg[6][8]  ( .D(\stage_1_output[6][8] ), .CP(clk), 
        .Q(\stage_1_retimer[6][8] ) );
  DFQD1 \stage_1_retimer_reg[6][7]  ( .D(\stage_1_output[6][7] ), .CP(clk), 
        .Q(\stage_1_retimer[6][7] ) );
  DFQD1 \stage_1_retimer_reg[6][6]  ( .D(\stage_1_output[6][6] ), .CP(clk), 
        .Q(\stage_1_retimer[6][6] ) );
  DFQD1 \stage_1_retimer_reg[6][5]  ( .D(\stage_1_output[6][5] ), .CP(clk), 
        .Q(\stage_1_retimer[6][5] ) );
  DFQD1 \stage_1_retimer_reg[6][4]  ( .D(\stage_1_output[6][4] ), .CP(clk), 
        .Q(\stage_1_retimer[6][4] ) );
  DFQD1 \stage_1_retimer_reg[6][3]  ( .D(\stage_1_output[6][3] ), .CP(clk), 
        .Q(\stage_1_retimer[6][3] ) );
  DFQD1 \stage_1_retimer_reg[6][2]  ( .D(\stage_1_output[6][2] ), .CP(clk), 
        .Q(\stage_1_retimer[6][2] ) );
  DFQD1 \stage_1_retimer_reg[6][1]  ( .D(\stage_1_output[6][1] ), .CP(clk), 
        .Q(\stage_1_retimer[6][1] ) );
  DFQD1 \stage_1_retimer_reg[6][0]  ( .D(\stage_1_output[6][0] ), .CP(clk), 
        .Q(\stage_1_retimer[6][0] ) );
  DFQD1 \stage_1_retimer_reg[5][19]  ( .D(\stage_1_output[5][19] ), .CP(clk), 
        .Q(\stage_1_retimer[5][19] ) );
  DFQD1 \stage_1_retimer_reg[5][18]  ( .D(\stage_1_output[5][18] ), .CP(clk), 
        .Q(\stage_1_retimer[5][18] ) );
  DFQD1 \stage_1_retimer_reg[5][17]  ( .D(\stage_1_output[5][17] ), .CP(clk), 
        .Q(\stage_1_retimer[5][17] ) );
  DFQD1 \stage_1_retimer_reg[5][16]  ( .D(\stage_1_output[5][16] ), .CP(clk), 
        .Q(\stage_1_retimer[5][16] ) );
  DFQD1 \stage_1_retimer_reg[5][15]  ( .D(\stage_1_output[5][15] ), .CP(clk), 
        .Q(\stage_1_retimer[5][15] ) );
  DFQD1 \stage_1_retimer_reg[5][14]  ( .D(\stage_1_output[5][14] ), .CP(clk), 
        .Q(\stage_1_retimer[5][14] ) );
  DFQD1 \stage_1_retimer_reg[5][13]  ( .D(\stage_1_output[5][13] ), .CP(clk), 
        .Q(\stage_1_retimer[5][13] ) );
  DFQD1 \stage_1_retimer_reg[5][12]  ( .D(\stage_1_output[5][12] ), .CP(clk), 
        .Q(\stage_1_retimer[5][12] ) );
  DFQD1 \stage_1_retimer_reg[5][11]  ( .D(\stage_1_output[5][11] ), .CP(clk), 
        .Q(\stage_1_retimer[5][11] ) );
  DFQD1 \stage_1_retimer_reg[5][10]  ( .D(\stage_1_output[5][10] ), .CP(clk), 
        .Q(\stage_1_retimer[5][10] ) );
  DFQD1 \stage_1_retimer_reg[5][9]  ( .D(\stage_1_output[5][9] ), .CP(clk), 
        .Q(\stage_1_retimer[5][9] ) );
  DFQD1 \stage_1_retimer_reg[5][8]  ( .D(\stage_1_output[5][8] ), .CP(clk), 
        .Q(\stage_1_retimer[5][8] ) );
  DFQD1 \stage_1_retimer_reg[5][7]  ( .D(\stage_1_output[5][7] ), .CP(clk), 
        .Q(\stage_1_retimer[5][7] ) );
  DFQD1 \stage_1_retimer_reg[5][6]  ( .D(\stage_1_output[5][6] ), .CP(clk), 
        .Q(\stage_1_retimer[5][6] ) );
  DFQD1 \stage_1_retimer_reg[5][5]  ( .D(\stage_1_output[5][5] ), .CP(clk), 
        .Q(\stage_1_retimer[5][5] ) );
  DFQD1 \stage_1_retimer_reg[5][4]  ( .D(\stage_1_output[5][4] ), .CP(clk), 
        .Q(\stage_1_retimer[5][4] ) );
  DFQD1 \stage_1_retimer_reg[5][3]  ( .D(\stage_1_output[5][3] ), .CP(clk), 
        .Q(\stage_1_retimer[5][3] ) );
  DFQD1 \stage_1_retimer_reg[5][2]  ( .D(\stage_1_output[5][2] ), .CP(clk), 
        .Q(\stage_1_retimer[5][2] ) );
  DFQD1 \stage_1_retimer_reg[5][1]  ( .D(\stage_1_output[5][1] ), .CP(clk), 
        .Q(\stage_1_retimer[5][1] ) );
  DFQD1 \stage_1_retimer_reg[5][0]  ( .D(\stage_1_output[5][0] ), .CP(clk), 
        .Q(\stage_1_retimer[5][0] ) );
  DFQD1 \stage_1_retimer_reg[4][19]  ( .D(\stage_1_output[4][19] ), .CP(clk), 
        .Q(\stage_1_retimer[4][19] ) );
  DFQD1 \stage_1_retimer_reg[4][18]  ( .D(\stage_1_output[4][18] ), .CP(clk), 
        .Q(\stage_1_retimer[4][18] ) );
  DFQD1 \stage_1_retimer_reg[4][17]  ( .D(\stage_1_output[4][17] ), .CP(clk), 
        .Q(\stage_1_retimer[4][17] ) );
  DFQD1 \stage_1_retimer_reg[4][16]  ( .D(\stage_1_output[4][16] ), .CP(clk), 
        .Q(\stage_1_retimer[4][16] ) );
  DFQD1 \stage_1_retimer_reg[4][15]  ( .D(\stage_1_output[4][15] ), .CP(clk), 
        .Q(\stage_1_retimer[4][15] ) );
  DFQD1 \stage_1_retimer_reg[4][14]  ( .D(\stage_1_output[4][14] ), .CP(clk), 
        .Q(\stage_1_retimer[4][14] ) );
  DFQD1 \stage_1_retimer_reg[4][13]  ( .D(\stage_1_output[4][13] ), .CP(clk), 
        .Q(\stage_1_retimer[4][13] ) );
  DFQD1 \stage_1_retimer_reg[4][12]  ( .D(\stage_1_output[4][12] ), .CP(clk), 
        .Q(\stage_1_retimer[4][12] ) );
  DFQD1 \stage_1_retimer_reg[4][11]  ( .D(\stage_1_output[4][11] ), .CP(clk), 
        .Q(\stage_1_retimer[4][11] ) );
  DFQD1 \stage_1_retimer_reg[4][10]  ( .D(\stage_1_output[4][10] ), .CP(clk), 
        .Q(\stage_1_retimer[4][10] ) );
  DFQD1 \stage_1_retimer_reg[4][9]  ( .D(\stage_1_output[4][9] ), .CP(clk), 
        .Q(\stage_1_retimer[4][9] ) );
  DFQD1 \stage_1_retimer_reg[4][8]  ( .D(\stage_1_output[4][8] ), .CP(clk), 
        .Q(\stage_1_retimer[4][8] ) );
  DFQD1 \stage_1_retimer_reg[4][7]  ( .D(\stage_1_output[4][7] ), .CP(clk), 
        .Q(\stage_1_retimer[4][7] ) );
  DFQD1 \stage_1_retimer_reg[4][6]  ( .D(\stage_1_output[4][6] ), .CP(clk), 
        .Q(\stage_1_retimer[4][6] ) );
  DFQD1 \stage_1_retimer_reg[4][5]  ( .D(\stage_1_output[4][5] ), .CP(clk), 
        .Q(\stage_1_retimer[4][5] ) );
  DFQD1 \stage_1_retimer_reg[4][4]  ( .D(\stage_1_output[4][4] ), .CP(clk), 
        .Q(\stage_1_retimer[4][4] ) );
  DFQD1 \stage_1_retimer_reg[4][3]  ( .D(\stage_1_output[4][3] ), .CP(clk), 
        .Q(\stage_1_retimer[4][3] ) );
  DFQD1 \stage_1_retimer_reg[4][2]  ( .D(\stage_1_output[4][2] ), .CP(clk), 
        .Q(\stage_1_retimer[4][2] ) );
  DFQD1 \stage_1_retimer_reg[4][1]  ( .D(\stage_1_output[4][1] ), .CP(clk), 
        .Q(\stage_1_retimer[4][1] ) );
  DFQD1 \stage_1_retimer_reg[4][0]  ( .D(\stage_1_output[4][0] ), .CP(clk), 
        .Q(\stage_1_retimer[4][0] ) );
  DFQD1 \stage_1_retimer_reg[3][19]  ( .D(\stage_1_output[3][19] ), .CP(clk), 
        .Q(\stage_1_retimer[3][19] ) );
  DFQD1 \stage_1_retimer_reg[3][18]  ( .D(\stage_1_output[3][18] ), .CP(clk), 
        .Q(\stage_1_retimer[3][18] ) );
  DFQD1 \stage_1_retimer_reg[3][17]  ( .D(\stage_1_output[3][17] ), .CP(clk), 
        .Q(\stage_1_retimer[3][17] ) );
  DFQD1 \stage_1_retimer_reg[3][16]  ( .D(\stage_1_output[3][16] ), .CP(clk), 
        .Q(\stage_1_retimer[3][16] ) );
  DFQD1 \stage_1_retimer_reg[3][15]  ( .D(\stage_1_output[3][15] ), .CP(clk), 
        .Q(\stage_1_retimer[3][15] ) );
  DFQD1 \stage_1_retimer_reg[3][14]  ( .D(\stage_1_output[3][14] ), .CP(clk), 
        .Q(\stage_1_retimer[3][14] ) );
  DFQD1 \stage_1_retimer_reg[3][13]  ( .D(\stage_1_output[3][13] ), .CP(clk), 
        .Q(\stage_1_retimer[3][13] ) );
  DFQD1 \stage_1_retimer_reg[3][12]  ( .D(\stage_1_output[3][12] ), .CP(clk), 
        .Q(\stage_1_retimer[3][12] ) );
  DFQD1 \stage_1_retimer_reg[3][11]  ( .D(\stage_1_output[3][11] ), .CP(clk), 
        .Q(\stage_1_retimer[3][11] ) );
  DFQD1 \stage_1_retimer_reg[3][10]  ( .D(\stage_1_output[3][10] ), .CP(clk), 
        .Q(\stage_1_retimer[3][10] ) );
  DFQD1 \stage_1_retimer_reg[3][9]  ( .D(\stage_1_output[3][9] ), .CP(clk), 
        .Q(\stage_1_retimer[3][9] ) );
  DFQD1 \stage_1_retimer_reg[3][8]  ( .D(\stage_1_output[3][8] ), .CP(clk), 
        .Q(\stage_1_retimer[3][8] ) );
  DFQD1 \stage_1_retimer_reg[3][7]  ( .D(\stage_1_output[3][7] ), .CP(clk), 
        .Q(\stage_1_retimer[3][7] ) );
  DFQD1 \stage_1_retimer_reg[3][6]  ( .D(\stage_1_output[3][6] ), .CP(clk), 
        .Q(\stage_1_retimer[3][6] ) );
  DFQD1 \stage_1_retimer_reg[3][5]  ( .D(\stage_1_output[3][5] ), .CP(clk), 
        .Q(\stage_1_retimer[3][5] ) );
  DFQD1 \stage_1_retimer_reg[3][4]  ( .D(\stage_1_output[3][4] ), .CP(clk), 
        .Q(\stage_1_retimer[3][4] ) );
  DFQD1 \stage_1_retimer_reg[3][3]  ( .D(\stage_1_output[3][3] ), .CP(clk), 
        .Q(\stage_1_retimer[3][3] ) );
  DFQD1 \stage_1_retimer_reg[3][2]  ( .D(\stage_1_output[3][2] ), .CP(clk), 
        .Q(\stage_1_retimer[3][2] ) );
  DFQD1 \stage_1_retimer_reg[3][1]  ( .D(\stage_1_output[3][1] ), .CP(clk), 
        .Q(\stage_1_retimer[3][1] ) );
  DFQD1 \stage_1_retimer_reg[3][0]  ( .D(\stage_1_output[3][0] ), .CP(clk), 
        .Q(\stage_1_retimer[3][0] ) );
  DFQD1 \stage_1_retimer_reg[2][19]  ( .D(\stage_1_output[2][19] ), .CP(clk), 
        .Q(\stage_1_retimer[2][19] ) );
  DFQD1 \stage_1_retimer_reg[2][18]  ( .D(\stage_1_output[2][18] ), .CP(clk), 
        .Q(\stage_1_retimer[2][18] ) );
  DFQD1 \stage_1_retimer_reg[2][17]  ( .D(\stage_1_output[2][17] ), .CP(clk), 
        .Q(\stage_1_retimer[2][17] ) );
  DFQD1 \stage_1_retimer_reg[2][16]  ( .D(\stage_1_output[2][16] ), .CP(clk), 
        .Q(\stage_1_retimer[2][16] ) );
  DFQD1 \stage_1_retimer_reg[2][15]  ( .D(\stage_1_output[2][15] ), .CP(clk), 
        .Q(\stage_1_retimer[2][15] ) );
  DFQD1 \stage_1_retimer_reg[2][14]  ( .D(\stage_1_output[2][14] ), .CP(clk), 
        .Q(\stage_1_retimer[2][14] ) );
  DFQD1 \stage_1_retimer_reg[2][13]  ( .D(\stage_1_output[2][13] ), .CP(clk), 
        .Q(\stage_1_retimer[2][13] ) );
  DFQD1 \stage_1_retimer_reg[2][12]  ( .D(\stage_1_output[2][12] ), .CP(clk), 
        .Q(\stage_1_retimer[2][12] ) );
  DFQD1 \stage_1_retimer_reg[2][11]  ( .D(\stage_1_output[2][11] ), .CP(clk), 
        .Q(\stage_1_retimer[2][11] ) );
  DFQD1 \stage_1_retimer_reg[2][10]  ( .D(\stage_1_output[2][10] ), .CP(clk), 
        .Q(\stage_1_retimer[2][10] ) );
  DFQD1 \stage_1_retimer_reg[2][9]  ( .D(\stage_1_output[2][9] ), .CP(clk), 
        .Q(\stage_1_retimer[2][9] ) );
  DFQD1 \stage_1_retimer_reg[2][8]  ( .D(\stage_1_output[2][8] ), .CP(clk), 
        .Q(\stage_1_retimer[2][8] ) );
  DFQD1 \stage_1_retimer_reg[2][7]  ( .D(\stage_1_output[2][7] ), .CP(clk), 
        .Q(\stage_1_retimer[2][7] ) );
  DFQD1 \stage_1_retimer_reg[2][6]  ( .D(\stage_1_output[2][6] ), .CP(clk), 
        .Q(\stage_1_retimer[2][6] ) );
  DFQD1 \stage_1_retimer_reg[2][5]  ( .D(\stage_1_output[2][5] ), .CP(clk), 
        .Q(\stage_1_retimer[2][5] ) );
  DFQD1 \stage_1_retimer_reg[2][4]  ( .D(\stage_1_output[2][4] ), .CP(clk), 
        .Q(\stage_1_retimer[2][4] ) );
  DFQD1 \stage_1_retimer_reg[2][3]  ( .D(\stage_1_output[2][3] ), .CP(clk), 
        .Q(\stage_1_retimer[2][3] ) );
  DFQD1 \stage_1_retimer_reg[2][2]  ( .D(\stage_1_output[2][2] ), .CP(clk), 
        .Q(\stage_1_retimer[2][2] ) );
  DFQD1 \stage_1_retimer_reg[2][1]  ( .D(\stage_1_output[2][1] ), .CP(clk), 
        .Q(\stage_1_retimer[2][1] ) );
  DFQD1 \stage_1_retimer_reg[2][0]  ( .D(\stage_1_output[2][0] ), .CP(clk), 
        .Q(\stage_1_retimer[2][0] ) );
  DFQD1 \stage_1_retimer_reg[1][19]  ( .D(\stage_1_output[1][19] ), .CP(clk), 
        .Q(\stage_1_retimer[1][19] ) );
  DFQD1 \stage_1_retimer_reg[1][18]  ( .D(\stage_1_output[1][18] ), .CP(clk), 
        .Q(\stage_1_retimer[1][18] ) );
  DFQD1 \stage_1_retimer_reg[1][17]  ( .D(\stage_1_output[1][17] ), .CP(clk), 
        .Q(\stage_1_retimer[1][17] ) );
  DFQD1 \stage_1_retimer_reg[1][16]  ( .D(\stage_1_output[1][16] ), .CP(clk), 
        .Q(\stage_1_retimer[1][16] ) );
  DFQD1 \stage_1_retimer_reg[1][15]  ( .D(\stage_1_output[1][15] ), .CP(clk), 
        .Q(\stage_1_retimer[1][15] ) );
  DFQD1 \stage_1_retimer_reg[1][14]  ( .D(\stage_1_output[1][14] ), .CP(clk), 
        .Q(\stage_1_retimer[1][14] ) );
  DFQD1 \stage_1_retimer_reg[1][13]  ( .D(\stage_1_output[1][13] ), .CP(clk), 
        .Q(\stage_1_retimer[1][13] ) );
  DFQD1 \stage_1_retimer_reg[1][12]  ( .D(\stage_1_output[1][12] ), .CP(clk), 
        .Q(\stage_1_retimer[1][12] ) );
  DFQD1 \stage_1_retimer_reg[1][11]  ( .D(\stage_1_output[1][11] ), .CP(clk), 
        .Q(\stage_1_retimer[1][11] ) );
  DFQD1 \stage_1_retimer_reg[1][10]  ( .D(\stage_1_output[1][10] ), .CP(clk), 
        .Q(\stage_1_retimer[1][10] ) );
  DFQD1 \stage_1_retimer_reg[1][9]  ( .D(\stage_1_output[1][9] ), .CP(clk), 
        .Q(\stage_1_retimer[1][9] ) );
  DFQD1 \stage_1_retimer_reg[1][8]  ( .D(\stage_1_output[1][8] ), .CP(clk), 
        .Q(\stage_1_retimer[1][8] ) );
  DFQD1 \stage_1_retimer_reg[1][7]  ( .D(\stage_1_output[1][7] ), .CP(clk), 
        .Q(\stage_1_retimer[1][7] ) );
  DFQD1 \stage_1_retimer_reg[1][6]  ( .D(\stage_1_output[1][6] ), .CP(clk), 
        .Q(\stage_1_retimer[1][6] ) );
  DFQD1 \stage_1_retimer_reg[1][5]  ( .D(\stage_1_output[1][5] ), .CP(clk), 
        .Q(\stage_1_retimer[1][5] ) );
  DFQD1 \stage_1_retimer_reg[1][4]  ( .D(\stage_1_output[1][4] ), .CP(clk), 
        .Q(\stage_1_retimer[1][4] ) );
  DFQD1 \stage_1_retimer_reg[1][3]  ( .D(\stage_1_output[1][3] ), .CP(clk), 
        .Q(\stage_1_retimer[1][3] ) );
  DFQD1 \stage_1_retimer_reg[1][2]  ( .D(\stage_1_output[1][2] ), .CP(clk), 
        .Q(\stage_1_retimer[1][2] ) );
  DFQD1 \stage_1_retimer_reg[1][1]  ( .D(\stage_1_output[1][1] ), .CP(clk), 
        .Q(\stage_1_retimer[1][1] ) );
  DFQD1 \stage_1_retimer_reg[1][0]  ( .D(\stage_1_output[1][0] ), .CP(clk), 
        .Q(\stage_1_retimer[1][0] ) );
  DFQD1 \stage_1_retimer_reg[0][19]  ( .D(\stage_1_output[0][19] ), .CP(clk), 
        .Q(\stage_1_retimer[0][19] ) );
  DFQD1 \stage_1_retimer_reg[0][18]  ( .D(\stage_1_output[0][18] ), .CP(clk), 
        .Q(\stage_1_retimer[0][18] ) );
  DFQD1 \stage_1_retimer_reg[0][17]  ( .D(\stage_1_output[0][17] ), .CP(clk), 
        .Q(\stage_1_retimer[0][17] ) );
  DFQD1 \stage_1_retimer_reg[0][16]  ( .D(\stage_1_output[0][16] ), .CP(clk), 
        .Q(\stage_1_retimer[0][16] ) );
  DFQD1 \stage_1_retimer_reg[0][15]  ( .D(\stage_1_output[0][15] ), .CP(clk), 
        .Q(\stage_1_retimer[0][15] ) );
  DFQD1 \stage_1_retimer_reg[0][14]  ( .D(\stage_1_output[0][14] ), .CP(clk), 
        .Q(\stage_1_retimer[0][14] ) );
  DFQD1 \stage_1_retimer_reg[0][13]  ( .D(\stage_1_output[0][13] ), .CP(clk), 
        .Q(\stage_1_retimer[0][13] ) );
  DFQD1 \stage_1_retimer_reg[0][12]  ( .D(\stage_1_output[0][12] ), .CP(clk), 
        .Q(\stage_1_retimer[0][12] ) );
  DFQD1 \stage_1_retimer_reg[0][11]  ( .D(\stage_1_output[0][11] ), .CP(clk), 
        .Q(\stage_1_retimer[0][11] ) );
  DFQD1 \stage_1_retimer_reg[0][10]  ( .D(\stage_1_output[0][10] ), .CP(clk), 
        .Q(\stage_1_retimer[0][10] ) );
  DFQD1 \stage_1_retimer_reg[0][9]  ( .D(\stage_1_output[0][9] ), .CP(clk), 
        .Q(\stage_1_retimer[0][9] ) );
  DFQD1 \stage_1_retimer_reg[0][8]  ( .D(\stage_1_output[0][8] ), .CP(clk), 
        .Q(\stage_1_retimer[0][8] ) );
  DFQD1 \stage_1_retimer_reg[0][7]  ( .D(\stage_1_output[0][7] ), .CP(clk), 
        .Q(\stage_1_retimer[0][7] ) );
  DFQD1 \stage_1_retimer_reg[0][6]  ( .D(\stage_1_output[0][6] ), .CP(clk), 
        .Q(\stage_1_retimer[0][6] ) );
  DFQD1 \stage_1_retimer_reg[0][5]  ( .D(\stage_1_output[0][5] ), .CP(clk), 
        .Q(\stage_1_retimer[0][5] ) );
  DFQD1 \stage_1_retimer_reg[0][4]  ( .D(\stage_1_output[0][4] ), .CP(clk), 
        .Q(\stage_1_retimer[0][4] ) );
  DFQD1 \stage_1_retimer_reg[0][3]  ( .D(\stage_1_output[0][3] ), .CP(clk), 
        .Q(\stage_1_retimer[0][3] ) );
  DFQD1 \stage_1_retimer_reg[0][2]  ( .D(\stage_1_output[0][2] ), .CP(clk), 
        .Q(\stage_1_retimer[0][2] ) );
  DFQD1 \stage_1_retimer_reg[0][1]  ( .D(\stage_1_output[0][1] ), .CP(clk), 
        .Q(\stage_1_retimer[0][1] ) );
  DFQD1 \stage_1_retimer_reg[0][0]  ( .D(\stage_1_output[0][0] ), .CP(clk), 
        .Q(\stage_1_retimer[0][0] ) );
  DFQD1 \stage_2_retimer_reg[7][19]  ( .D(\stage_2_output[7][19] ), .CP(clk), 
        .Q(\stage_2_retimer[7][19] ) );
  DFQD1 \stage_2_retimer_reg[7][18]  ( .D(\stage_2_output[7][18] ), .CP(clk), 
        .Q(\stage_2_retimer[7][18] ) );
  DFQD1 \stage_2_retimer_reg[7][17]  ( .D(\stage_2_output[7][17] ), .CP(clk), 
        .Q(\stage_2_retimer[7][17] ) );
  DFQD1 \stage_2_retimer_reg[7][16]  ( .D(\stage_2_output[7][16] ), .CP(clk), 
        .Q(\stage_2_retimer[7][16] ) );
  DFQD1 \stage_2_retimer_reg[7][15]  ( .D(\stage_2_output[7][15] ), .CP(clk), 
        .Q(\stage_2_retimer[7][15] ) );
  DFQD1 \stage_2_retimer_reg[7][14]  ( .D(\stage_2_output[7][14] ), .CP(clk), 
        .Q(\stage_2_retimer[7][14] ) );
  DFQD1 \stage_2_retimer_reg[7][13]  ( .D(\stage_2_output[7][13] ), .CP(clk), 
        .Q(\stage_2_retimer[7][13] ) );
  DFQD1 \stage_2_retimer_reg[7][12]  ( .D(\stage_2_output[7][12] ), .CP(clk), 
        .Q(\stage_2_retimer[7][12] ) );
  DFQD1 \stage_2_retimer_reg[7][11]  ( .D(\stage_2_output[7][11] ), .CP(clk), 
        .Q(\stage_2_retimer[7][11] ) );
  DFQD1 \stage_2_retimer_reg[7][10]  ( .D(\stage_2_output[7][10] ), .CP(clk), 
        .Q(\stage_2_retimer[7][10] ) );
  DFQD1 \stage_2_retimer_reg[7][9]  ( .D(\stage_2_output[7][9] ), .CP(clk), 
        .Q(\stage_2_retimer[7][9] ) );
  DFQD1 \stage_2_retimer_reg[7][8]  ( .D(\stage_2_output[7][8] ), .CP(clk), 
        .Q(\stage_2_retimer[7][8] ) );
  DFQD1 \stage_2_retimer_reg[7][7]  ( .D(\stage_2_output[7][7] ), .CP(clk), 
        .Q(\stage_2_retimer[7][7] ) );
  DFQD1 \stage_2_retimer_reg[7][6]  ( .D(\stage_2_output[7][6] ), .CP(clk), 
        .Q(\stage_2_retimer[7][6] ) );
  DFQD1 \stage_2_retimer_reg[7][5]  ( .D(\stage_2_output[7][5] ), .CP(clk), 
        .Q(\stage_2_retimer[7][5] ) );
  DFQD1 \stage_2_retimer_reg[7][4]  ( .D(\stage_2_output[7][4] ), .CP(clk), 
        .Q(\stage_2_retimer[7][4] ) );
  DFQD1 \stage_2_retimer_reg[7][3]  ( .D(\stage_2_output[7][3] ), .CP(clk), 
        .Q(\stage_2_retimer[7][3] ) );
  DFQD1 \stage_2_retimer_reg[7][2]  ( .D(\stage_2_output[7][2] ), .CP(clk), 
        .Q(\stage_2_retimer[7][2] ) );
  DFQD1 \stage_2_retimer_reg[7][1]  ( .D(\stage_2_output[7][1] ), .CP(clk), 
        .Q(\stage_2_retimer[7][1] ) );
  DFQD1 \stage_2_retimer_reg[7][0]  ( .D(\stage_2_output[7][0] ), .CP(clk), 
        .Q(\stage_2_retimer[7][0] ) );
  DFQD1 \stage_2_retimer_reg[6][19]  ( .D(\stage_2_output[6][19] ), .CP(clk), 
        .Q(\stage_2_retimer[6][19] ) );
  DFQD1 \stage_2_retimer_reg[6][18]  ( .D(\stage_2_output[6][18] ), .CP(clk), 
        .Q(\stage_2_retimer[6][18] ) );
  DFQD1 \stage_2_retimer_reg[6][17]  ( .D(\stage_2_output[6][17] ), .CP(clk), 
        .Q(\stage_2_retimer[6][17] ) );
  DFQD1 \stage_2_retimer_reg[6][16]  ( .D(\stage_2_output[6][16] ), .CP(clk), 
        .Q(\stage_2_retimer[6][16] ) );
  DFQD1 \stage_2_retimer_reg[6][15]  ( .D(\stage_2_output[6][15] ), .CP(clk), 
        .Q(\stage_2_retimer[6][15] ) );
  DFQD1 \stage_2_retimer_reg[6][14]  ( .D(\stage_2_output[6][14] ), .CP(clk), 
        .Q(\stage_2_retimer[6][14] ) );
  DFQD1 \stage_2_retimer_reg[6][13]  ( .D(\stage_2_output[6][13] ), .CP(clk), 
        .Q(\stage_2_retimer[6][13] ) );
  DFQD1 \stage_2_retimer_reg[6][12]  ( .D(\stage_2_output[6][12] ), .CP(clk), 
        .Q(\stage_2_retimer[6][12] ) );
  DFQD1 \stage_2_retimer_reg[6][11]  ( .D(\stage_2_output[6][11] ), .CP(clk), 
        .Q(\stage_2_retimer[6][11] ) );
  DFQD1 \stage_2_retimer_reg[6][10]  ( .D(\stage_2_output[6][10] ), .CP(clk), 
        .Q(\stage_2_retimer[6][10] ) );
  DFQD1 \stage_2_retimer_reg[6][9]  ( .D(\stage_2_output[6][9] ), .CP(clk), 
        .Q(\stage_2_retimer[6][9] ) );
  DFQD1 \stage_2_retimer_reg[6][8]  ( .D(\stage_2_output[6][8] ), .CP(clk), 
        .Q(\stage_2_retimer[6][8] ) );
  DFQD1 \stage_2_retimer_reg[6][7]  ( .D(\stage_2_output[6][7] ), .CP(clk), 
        .Q(\stage_2_retimer[6][7] ) );
  DFQD1 \stage_2_retimer_reg[6][6]  ( .D(\stage_2_output[6][6] ), .CP(clk), 
        .Q(\stage_2_retimer[6][6] ) );
  DFQD1 \stage_2_retimer_reg[6][5]  ( .D(\stage_2_output[6][5] ), .CP(clk), 
        .Q(\stage_2_retimer[6][5] ) );
  DFQD1 \stage_2_retimer_reg[6][4]  ( .D(\stage_2_output[6][4] ), .CP(clk), 
        .Q(\stage_2_retimer[6][4] ) );
  DFQD1 \stage_2_retimer_reg[6][3]  ( .D(\stage_2_output[6][3] ), .CP(clk), 
        .Q(\stage_2_retimer[6][3] ) );
  DFQD1 \stage_2_retimer_reg[6][2]  ( .D(\stage_2_output[6][2] ), .CP(clk), 
        .Q(\stage_2_retimer[6][2] ) );
  DFQD1 \stage_2_retimer_reg[6][1]  ( .D(\stage_2_output[6][1] ), .CP(clk), 
        .Q(\stage_2_retimer[6][1] ) );
  DFQD1 \stage_2_retimer_reg[6][0]  ( .D(\stage_2_output[6][0] ), .CP(clk), 
        .Q(\stage_2_retimer[6][0] ) );
  DFQD1 \stage_2_retimer_reg[5][19]  ( .D(\stage_2_output[5][19] ), .CP(clk), 
        .Q(\stage_2_retimer[5][19] ) );
  DFQD1 \stage_2_retimer_reg[5][18]  ( .D(\stage_2_output[5][18] ), .CP(clk), 
        .Q(\stage_2_retimer[5][18] ) );
  DFQD1 \stage_2_retimer_reg[5][17]  ( .D(\stage_2_output[5][17] ), .CP(clk), 
        .Q(\stage_2_retimer[5][17] ) );
  DFQD1 \stage_2_retimer_reg[5][16]  ( .D(\stage_2_output[5][16] ), .CP(clk), 
        .Q(\stage_2_retimer[5][16] ) );
  DFQD1 \stage_2_retimer_reg[5][15]  ( .D(\stage_2_output[5][15] ), .CP(clk), 
        .Q(\stage_2_retimer[5][15] ) );
  DFQD1 \stage_2_retimer_reg[5][14]  ( .D(\stage_2_output[5][14] ), .CP(clk), 
        .Q(\stage_2_retimer[5][14] ) );
  DFQD1 \stage_2_retimer_reg[5][13]  ( .D(\stage_2_output[5][13] ), .CP(clk), 
        .Q(\stage_2_retimer[5][13] ) );
  DFQD1 \stage_2_retimer_reg[5][12]  ( .D(\stage_2_output[5][12] ), .CP(clk), 
        .Q(\stage_2_retimer[5][12] ) );
  DFQD1 \stage_2_retimer_reg[5][11]  ( .D(\stage_2_output[5][11] ), .CP(clk), 
        .Q(\stage_2_retimer[5][11] ) );
  DFQD1 \stage_2_retimer_reg[5][10]  ( .D(\stage_2_output[5][10] ), .CP(clk), 
        .Q(\stage_2_retimer[5][10] ) );
  DFQD1 \stage_2_retimer_reg[5][9]  ( .D(\stage_2_output[5][9] ), .CP(clk), 
        .Q(\stage_2_retimer[5][9] ) );
  DFQD1 \stage_2_retimer_reg[5][8]  ( .D(\stage_2_output[5][8] ), .CP(clk), 
        .Q(\stage_2_retimer[5][8] ) );
  DFQD1 \stage_2_retimer_reg[5][7]  ( .D(\stage_2_output[5][7] ), .CP(clk), 
        .Q(\stage_2_retimer[5][7] ) );
  DFQD1 \stage_2_retimer_reg[5][6]  ( .D(\stage_2_output[5][6] ), .CP(clk), 
        .Q(\stage_2_retimer[5][6] ) );
  DFQD1 \stage_2_retimer_reg[5][5]  ( .D(\stage_2_output[5][5] ), .CP(clk), 
        .Q(\stage_2_retimer[5][5] ) );
  DFQD1 \stage_2_retimer_reg[5][4]  ( .D(\stage_2_output[5][4] ), .CP(clk), 
        .Q(\stage_2_retimer[5][4] ) );
  DFQD1 \stage_2_retimer_reg[5][3]  ( .D(\stage_2_output[5][3] ), .CP(clk), 
        .Q(\stage_2_retimer[5][3] ) );
  DFQD1 \stage_2_retimer_reg[5][2]  ( .D(\stage_2_output[5][2] ), .CP(clk), 
        .Q(\stage_2_retimer[5][2] ) );
  DFQD1 \stage_2_retimer_reg[5][1]  ( .D(\stage_2_output[5][1] ), .CP(clk), 
        .Q(\stage_2_retimer[5][1] ) );
  DFQD1 \stage_2_retimer_reg[5][0]  ( .D(\stage_2_output[5][0] ), .CP(clk), 
        .Q(\stage_2_retimer[5][0] ) );
  DFQD1 \stage_2_retimer_reg[4][19]  ( .D(\stage_2_output[4][19] ), .CP(clk), 
        .Q(\stage_2_retimer[4][19] ) );
  DFQD1 \stage_2_retimer_reg[4][18]  ( .D(\stage_2_output[4][18] ), .CP(clk), 
        .Q(\stage_2_retimer[4][18] ) );
  DFQD1 \stage_2_retimer_reg[4][17]  ( .D(\stage_2_output[4][17] ), .CP(clk), 
        .Q(\stage_2_retimer[4][17] ) );
  DFQD1 \stage_2_retimer_reg[4][16]  ( .D(\stage_2_output[4][16] ), .CP(clk), 
        .Q(\stage_2_retimer[4][16] ) );
  DFQD1 \stage_2_retimer_reg[4][15]  ( .D(\stage_2_output[4][15] ), .CP(clk), 
        .Q(\stage_2_retimer[4][15] ) );
  DFQD1 \stage_2_retimer_reg[4][14]  ( .D(\stage_2_output[4][14] ), .CP(clk), 
        .Q(\stage_2_retimer[4][14] ) );
  DFQD1 \stage_2_retimer_reg[4][13]  ( .D(\stage_2_output[4][13] ), .CP(clk), 
        .Q(\stage_2_retimer[4][13] ) );
  DFQD1 \stage_2_retimer_reg[4][12]  ( .D(\stage_2_output[4][12] ), .CP(clk), 
        .Q(\stage_2_retimer[4][12] ) );
  DFQD1 \stage_2_retimer_reg[4][11]  ( .D(\stage_2_output[4][11] ), .CP(clk), 
        .Q(\stage_2_retimer[4][11] ) );
  DFQD1 \stage_2_retimer_reg[4][10]  ( .D(\stage_2_output[4][10] ), .CP(clk), 
        .Q(\stage_2_retimer[4][10] ) );
  DFQD1 \stage_2_retimer_reg[4][9]  ( .D(\stage_2_output[4][9] ), .CP(clk), 
        .Q(\stage_2_retimer[4][9] ) );
  DFQD1 \stage_2_retimer_reg[4][8]  ( .D(\stage_2_output[4][8] ), .CP(clk), 
        .Q(\stage_2_retimer[4][8] ) );
  DFQD1 \stage_2_retimer_reg[4][7]  ( .D(\stage_2_output[4][7] ), .CP(clk), 
        .Q(\stage_2_retimer[4][7] ) );
  DFQD1 \stage_2_retimer_reg[4][6]  ( .D(\stage_2_output[4][6] ), .CP(clk), 
        .Q(\stage_2_retimer[4][6] ) );
  DFQD1 \stage_2_retimer_reg[4][5]  ( .D(\stage_2_output[4][5] ), .CP(clk), 
        .Q(\stage_2_retimer[4][5] ) );
  DFQD1 \stage_2_retimer_reg[4][4]  ( .D(\stage_2_output[4][4] ), .CP(clk), 
        .Q(\stage_2_retimer[4][4] ) );
  DFQD1 \stage_2_retimer_reg[4][3]  ( .D(\stage_2_output[4][3] ), .CP(clk), 
        .Q(\stage_2_retimer[4][3] ) );
  DFQD1 \stage_2_retimer_reg[4][2]  ( .D(\stage_2_output[4][2] ), .CP(clk), 
        .Q(\stage_2_retimer[4][2] ) );
  DFQD1 \stage_2_retimer_reg[4][1]  ( .D(\stage_2_output[4][1] ), .CP(clk), 
        .Q(\stage_2_retimer[4][1] ) );
  DFQD1 \stage_2_retimer_reg[4][0]  ( .D(\stage_2_output[4][0] ), .CP(clk), 
        .Q(\stage_2_retimer[4][0] ) );
  DFQD1 \stage_2_retimer_reg[3][19]  ( .D(\stage_2_output[3][19] ), .CP(clk), 
        .Q(\stage_2_retimer[3][19] ) );
  DFQD1 \stage_2_retimer_reg[3][18]  ( .D(\stage_2_output[3][18] ), .CP(clk), 
        .Q(\stage_2_retimer[3][18] ) );
  DFQD1 \stage_2_retimer_reg[3][17]  ( .D(\stage_2_output[3][17] ), .CP(clk), 
        .Q(\stage_2_retimer[3][17] ) );
  DFQD1 \stage_2_retimer_reg[3][16]  ( .D(\stage_2_output[3][16] ), .CP(clk), 
        .Q(\stage_2_retimer[3][16] ) );
  DFQD1 \stage_2_retimer_reg[3][15]  ( .D(\stage_2_output[3][15] ), .CP(clk), 
        .Q(\stage_2_retimer[3][15] ) );
  DFQD1 \stage_2_retimer_reg[3][14]  ( .D(\stage_2_output[3][14] ), .CP(clk), 
        .Q(\stage_2_retimer[3][14] ) );
  DFQD1 \stage_2_retimer_reg[3][13]  ( .D(\stage_2_output[3][13] ), .CP(clk), 
        .Q(\stage_2_retimer[3][13] ) );
  DFQD1 \stage_2_retimer_reg[3][12]  ( .D(\stage_2_output[3][12] ), .CP(clk), 
        .Q(\stage_2_retimer[3][12] ) );
  DFQD1 \stage_2_retimer_reg[3][11]  ( .D(\stage_2_output[3][11] ), .CP(clk), 
        .Q(\stage_2_retimer[3][11] ) );
  DFQD1 \stage_2_retimer_reg[3][10]  ( .D(\stage_2_output[3][10] ), .CP(clk), 
        .Q(\stage_2_retimer[3][10] ) );
  DFQD1 \stage_2_retimer_reg[3][9]  ( .D(\stage_2_output[3][9] ), .CP(clk), 
        .Q(\stage_2_retimer[3][9] ) );
  DFQD1 \stage_2_retimer_reg[3][8]  ( .D(\stage_2_output[3][8] ), .CP(clk), 
        .Q(\stage_2_retimer[3][8] ) );
  DFQD1 \stage_2_retimer_reg[3][7]  ( .D(\stage_2_output[3][7] ), .CP(clk), 
        .Q(\stage_2_retimer[3][7] ) );
  DFQD1 \stage_2_retimer_reg[3][6]  ( .D(\stage_2_output[3][6] ), .CP(clk), 
        .Q(\stage_2_retimer[3][6] ) );
  DFQD1 \stage_2_retimer_reg[3][5]  ( .D(\stage_2_output[3][5] ), .CP(clk), 
        .Q(\stage_2_retimer[3][5] ) );
  DFQD1 \stage_2_retimer_reg[3][4]  ( .D(\stage_2_output[3][4] ), .CP(clk), 
        .Q(\stage_2_retimer[3][4] ) );
  DFQD1 \stage_2_retimer_reg[3][3]  ( .D(\stage_2_output[3][3] ), .CP(clk), 
        .Q(\stage_2_retimer[3][3] ) );
  DFQD1 \stage_2_retimer_reg[3][2]  ( .D(\stage_2_output[3][2] ), .CP(clk), 
        .Q(\stage_2_retimer[3][2] ) );
  DFQD1 \stage_2_retimer_reg[3][1]  ( .D(\stage_2_output[3][1] ), .CP(clk), 
        .Q(\stage_2_retimer[3][1] ) );
  DFQD1 \stage_2_retimer_reg[3][0]  ( .D(\stage_2_output[3][0] ), .CP(clk), 
        .Q(\stage_2_retimer[3][0] ) );
  DFQD1 \stage_2_retimer_reg[2][19]  ( .D(\stage_2_output[2][19] ), .CP(clk), 
        .Q(\stage_2_retimer[2][19] ) );
  DFQD1 \stage_2_retimer_reg[2][18]  ( .D(\stage_2_output[2][18] ), .CP(clk), 
        .Q(\stage_2_retimer[2][18] ) );
  DFQD1 \stage_2_retimer_reg[2][17]  ( .D(\stage_2_output[2][17] ), .CP(clk), 
        .Q(\stage_2_retimer[2][17] ) );
  DFQD1 \stage_2_retimer_reg[2][16]  ( .D(\stage_2_output[2][16] ), .CP(clk), 
        .Q(\stage_2_retimer[2][16] ) );
  DFQD1 \stage_2_retimer_reg[2][15]  ( .D(\stage_2_output[2][15] ), .CP(clk), 
        .Q(\stage_2_retimer[2][15] ) );
  DFQD1 \stage_2_retimer_reg[2][14]  ( .D(\stage_2_output[2][14] ), .CP(clk), 
        .Q(\stage_2_retimer[2][14] ) );
  DFQD1 \stage_2_retimer_reg[2][13]  ( .D(\stage_2_output[2][13] ), .CP(clk), 
        .Q(\stage_2_retimer[2][13] ) );
  DFQD1 \stage_2_retimer_reg[2][12]  ( .D(\stage_2_output[2][12] ), .CP(clk), 
        .Q(\stage_2_retimer[2][12] ) );
  DFQD1 \stage_2_retimer_reg[2][11]  ( .D(\stage_2_output[2][11] ), .CP(clk), 
        .Q(\stage_2_retimer[2][11] ) );
  DFQD1 \stage_2_retimer_reg[2][10]  ( .D(\stage_2_output[2][10] ), .CP(clk), 
        .Q(\stage_2_retimer[2][10] ) );
  DFQD1 \stage_2_retimer_reg[2][9]  ( .D(\stage_2_output[2][9] ), .CP(clk), 
        .Q(\stage_2_retimer[2][9] ) );
  DFQD1 \stage_2_retimer_reg[2][8]  ( .D(\stage_2_output[2][8] ), .CP(clk), 
        .Q(\stage_2_retimer[2][8] ) );
  DFQD1 \stage_2_retimer_reg[2][7]  ( .D(\stage_2_output[2][7] ), .CP(clk), 
        .Q(\stage_2_retimer[2][7] ) );
  DFQD1 \stage_2_retimer_reg[2][6]  ( .D(\stage_2_output[2][6] ), .CP(clk), 
        .Q(\stage_2_retimer[2][6] ) );
  DFQD1 \stage_2_retimer_reg[2][5]  ( .D(\stage_2_output[2][5] ), .CP(clk), 
        .Q(\stage_2_retimer[2][5] ) );
  DFQD1 \stage_2_retimer_reg[2][4]  ( .D(\stage_2_output[2][4] ), .CP(clk), 
        .Q(\stage_2_retimer[2][4] ) );
  DFQD1 \stage_2_retimer_reg[2][3]  ( .D(\stage_2_output[2][3] ), .CP(clk), 
        .Q(\stage_2_retimer[2][3] ) );
  DFQD1 \stage_2_retimer_reg[2][2]  ( .D(\stage_2_output[2][2] ), .CP(clk), 
        .Q(\stage_2_retimer[2][2] ) );
  DFQD1 \stage_2_retimer_reg[2][1]  ( .D(\stage_2_output[2][1] ), .CP(clk), 
        .Q(\stage_2_retimer[2][1] ) );
  DFQD1 \stage_2_retimer_reg[2][0]  ( .D(\stage_2_output[2][0] ), .CP(clk), 
        .Q(\stage_2_retimer[2][0] ) );
  DFQD1 \stage_2_retimer_reg[1][19]  ( .D(\stage_2_output[1][19] ), .CP(clk), 
        .Q(\stage_2_retimer[1][19] ) );
  DFQD1 \stage_2_retimer_reg[1][18]  ( .D(\stage_2_output[1][18] ), .CP(clk), 
        .Q(\stage_2_retimer[1][18] ) );
  DFQD1 \stage_2_retimer_reg[1][17]  ( .D(\stage_2_output[1][17] ), .CP(clk), 
        .Q(\stage_2_retimer[1][17] ) );
  DFQD1 \stage_2_retimer_reg[1][16]  ( .D(\stage_2_output[1][16] ), .CP(clk), 
        .Q(\stage_2_retimer[1][16] ) );
  DFQD1 \stage_2_retimer_reg[1][15]  ( .D(\stage_2_output[1][15] ), .CP(clk), 
        .Q(\stage_2_retimer[1][15] ) );
  DFQD1 \stage_2_retimer_reg[1][14]  ( .D(\stage_2_output[1][14] ), .CP(clk), 
        .Q(\stage_2_retimer[1][14] ) );
  DFQD1 \stage_2_retimer_reg[1][13]  ( .D(\stage_2_output[1][13] ), .CP(clk), 
        .Q(\stage_2_retimer[1][13] ) );
  DFQD1 \stage_2_retimer_reg[1][12]  ( .D(\stage_2_output[1][12] ), .CP(clk), 
        .Q(\stage_2_retimer[1][12] ) );
  DFQD1 \stage_2_retimer_reg[1][11]  ( .D(\stage_2_output[1][11] ), .CP(clk), 
        .Q(\stage_2_retimer[1][11] ) );
  DFQD1 \stage_2_retimer_reg[1][10]  ( .D(\stage_2_output[1][10] ), .CP(clk), 
        .Q(\stage_2_retimer[1][10] ) );
  DFQD1 \stage_2_retimer_reg[1][9]  ( .D(\stage_2_output[1][9] ), .CP(clk), 
        .Q(\stage_2_retimer[1][9] ) );
  DFQD1 \stage_2_retimer_reg[1][8]  ( .D(\stage_2_output[1][8] ), .CP(clk), 
        .Q(\stage_2_retimer[1][8] ) );
  DFQD1 \stage_2_retimer_reg[1][7]  ( .D(\stage_2_output[1][7] ), .CP(clk), 
        .Q(\stage_2_retimer[1][7] ) );
  DFQD1 \stage_2_retimer_reg[1][6]  ( .D(\stage_2_output[1][6] ), .CP(clk), 
        .Q(\stage_2_retimer[1][6] ) );
  DFQD1 \stage_2_retimer_reg[1][5]  ( .D(\stage_2_output[1][5] ), .CP(clk), 
        .Q(\stage_2_retimer[1][5] ) );
  DFQD1 \stage_2_retimer_reg[1][4]  ( .D(\stage_2_output[1][4] ), .CP(clk), 
        .Q(\stage_2_retimer[1][4] ) );
  DFQD1 \stage_2_retimer_reg[1][3]  ( .D(\stage_2_output[1][3] ), .CP(clk), 
        .Q(\stage_2_retimer[1][3] ) );
  DFQD1 \stage_2_retimer_reg[1][2]  ( .D(\stage_2_output[1][2] ), .CP(clk), 
        .Q(\stage_2_retimer[1][2] ) );
  DFQD1 \stage_2_retimer_reg[1][1]  ( .D(\stage_2_output[1][1] ), .CP(clk), 
        .Q(\stage_2_retimer[1][1] ) );
  DFQD1 \stage_2_retimer_reg[1][0]  ( .D(\stage_2_output[1][0] ), .CP(clk), 
        .Q(\stage_2_retimer[1][0] ) );
  DFQD1 \stage_2_retimer_reg[0][19]  ( .D(\stage_2_output[0][19] ), .CP(clk), 
        .Q(\stage_2_retimer[0][19] ) );
  DFQD1 \stage_2_retimer_reg[0][18]  ( .D(\stage_2_output[0][18] ), .CP(clk), 
        .Q(\stage_2_retimer[0][18] ) );
  DFQD1 \stage_2_retimer_reg[0][17]  ( .D(\stage_2_output[0][17] ), .CP(clk), 
        .Q(\stage_2_retimer[0][17] ) );
  DFQD1 \stage_2_retimer_reg[0][16]  ( .D(\stage_2_output[0][16] ), .CP(clk), 
        .Q(\stage_2_retimer[0][16] ) );
  DFQD1 \stage_2_retimer_reg[0][15]  ( .D(\stage_2_output[0][15] ), .CP(clk), 
        .Q(\stage_2_retimer[0][15] ) );
  DFQD1 \stage_2_retimer_reg[0][14]  ( .D(\stage_2_output[0][14] ), .CP(clk), 
        .Q(\stage_2_retimer[0][14] ) );
  DFQD1 \stage_2_retimer_reg[0][13]  ( .D(\stage_2_output[0][13] ), .CP(clk), 
        .Q(\stage_2_retimer[0][13] ) );
  DFQD1 \stage_2_retimer_reg[0][12]  ( .D(\stage_2_output[0][12] ), .CP(clk), 
        .Q(\stage_2_retimer[0][12] ) );
  DFQD1 \stage_2_retimer_reg[0][11]  ( .D(\stage_2_output[0][11] ), .CP(clk), 
        .Q(\stage_2_retimer[0][11] ) );
  DFQD1 \stage_2_retimer_reg[0][10]  ( .D(\stage_2_output[0][10] ), .CP(clk), 
        .Q(\stage_2_retimer[0][10] ) );
  DFQD1 \stage_2_retimer_reg[0][9]  ( .D(\stage_2_output[0][9] ), .CP(clk), 
        .Q(\stage_2_retimer[0][9] ) );
  DFQD1 \stage_2_retimer_reg[0][8]  ( .D(\stage_2_output[0][8] ), .CP(clk), 
        .Q(\stage_2_retimer[0][8] ) );
  DFQD1 \stage_2_retimer_reg[0][7]  ( .D(\stage_2_output[0][7] ), .CP(clk), 
        .Q(\stage_2_retimer[0][7] ) );
  DFQD1 \stage_2_retimer_reg[0][6]  ( .D(\stage_2_output[0][6] ), .CP(clk), 
        .Q(\stage_2_retimer[0][6] ) );
  DFQD1 \stage_2_retimer_reg[0][5]  ( .D(\stage_2_output[0][5] ), .CP(clk), 
        .Q(\stage_2_retimer[0][5] ) );
  DFQD1 \stage_2_retimer_reg[0][4]  ( .D(\stage_2_output[0][4] ), .CP(clk), 
        .Q(\stage_2_retimer[0][4] ) );
  DFQD1 \stage_2_retimer_reg[0][3]  ( .D(\stage_2_output[0][3] ), .CP(clk), 
        .Q(\stage_2_retimer[0][3] ) );
  DFQD1 \stage_2_retimer_reg[0][2]  ( .D(\stage_2_output[0][2] ), .CP(clk), 
        .Q(\stage_2_retimer[0][2] ) );
  DFQD1 \stage_2_retimer_reg[0][1]  ( .D(\stage_2_output[0][1] ), .CP(clk), 
        .Q(\stage_2_retimer[0][1] ) );
  DFQD1 \stage_2_retimer_reg[0][0]  ( .D(\stage_2_output[0][0] ), .CP(clk), 
        .Q(\stage_2_retimer[0][0] ) );
  DFQD1 \stage_3_retimer_reg[7][19]  ( .D(\stage_3_output[7][19] ), .CP(clk), 
        .Q(\stage_3_retimer[7][19] ) );
  DFQD1 \stage_3_retimer_reg[7][18]  ( .D(\stage_3_output[7][18] ), .CP(clk), 
        .Q(\stage_3_retimer[7][18] ) );
  DFQD1 \stage_3_retimer_reg[7][17]  ( .D(\stage_3_output[7][17] ), .CP(clk), 
        .Q(\stage_3_retimer[7][17] ) );
  DFQD1 \stage_3_retimer_reg[7][16]  ( .D(\stage_3_output[7][16] ), .CP(clk), 
        .Q(\stage_3_retimer[7][16] ) );
  DFQD1 \stage_3_retimer_reg[7][15]  ( .D(\stage_3_output[7][15] ), .CP(clk), 
        .Q(\stage_3_retimer[7][15] ) );
  DFQD1 \stage_3_retimer_reg[7][14]  ( .D(\stage_3_output[7][14] ), .CP(clk), 
        .Q(\stage_3_retimer[7][14] ) );
  DFQD1 \stage_3_retimer_reg[7][13]  ( .D(\stage_3_output[7][13] ), .CP(clk), 
        .Q(\stage_3_retimer[7][13] ) );
  DFQD1 \stage_3_retimer_reg[7][12]  ( .D(\stage_3_output[7][12] ), .CP(clk), 
        .Q(\stage_3_retimer[7][12] ) );
  DFQD1 \stage_3_retimer_reg[7][11]  ( .D(\stage_3_output[7][11] ), .CP(clk), 
        .Q(\stage_3_retimer[7][11] ) );
  DFQD1 \stage_3_retimer_reg[7][10]  ( .D(\stage_3_output[7][10] ), .CP(clk), 
        .Q(\stage_3_retimer[7][10] ) );
  DFQD1 \stage_3_retimer_reg[7][9]  ( .D(\stage_3_output[7][9] ), .CP(clk), 
        .Q(\stage_3_retimer[7][9] ) );
  DFQD1 \stage_3_retimer_reg[7][8]  ( .D(\stage_3_output[7][8] ), .CP(clk), 
        .Q(\stage_3_retimer[7][8] ) );
  DFQD1 \stage_3_retimer_reg[7][7]  ( .D(\stage_3_output[7][7] ), .CP(clk), 
        .Q(\stage_3_retimer[7][7] ) );
  DFQD1 \stage_3_retimer_reg[7][6]  ( .D(\stage_3_output[7][6] ), .CP(clk), 
        .Q(\stage_3_retimer[7][6] ) );
  DFQD1 \stage_3_retimer_reg[7][5]  ( .D(\stage_3_output[7][5] ), .CP(clk), 
        .Q(\stage_3_retimer[7][5] ) );
  DFQD1 \stage_3_retimer_reg[7][4]  ( .D(\stage_3_output[7][4] ), .CP(clk), 
        .Q(\stage_3_retimer[7][4] ) );
  DFQD1 \stage_3_retimer_reg[7][3]  ( .D(\stage_3_output[7][3] ), .CP(clk), 
        .Q(\stage_3_retimer[7][3] ) );
  DFQD1 \stage_3_retimer_reg[7][2]  ( .D(\stage_3_output[7][2] ), .CP(clk), 
        .Q(\stage_3_retimer[7][2] ) );
  DFQD1 \stage_3_retimer_reg[7][1]  ( .D(\stage_3_output[7][1] ), .CP(clk), 
        .Q(\stage_3_retimer[7][1] ) );
  DFQD1 \stage_3_retimer_reg[7][0]  ( .D(\stage_3_output[7][0] ), .CP(clk), 
        .Q(\stage_3_retimer[7][0] ) );
  DFQD1 \stage_3_retimer_reg[6][19]  ( .D(\stage_3_output[6][19] ), .CP(clk), 
        .Q(\stage_3_retimer[6][19] ) );
  DFQD1 \stage_3_retimer_reg[6][18]  ( .D(\stage_3_output[6][18] ), .CP(clk), 
        .Q(\stage_3_retimer[6][18] ) );
  DFQD1 \stage_3_retimer_reg[6][17]  ( .D(\stage_3_output[6][17] ), .CP(clk), 
        .Q(\stage_3_retimer[6][17] ) );
  DFQD1 \stage_3_retimer_reg[6][16]  ( .D(\stage_3_output[6][16] ), .CP(clk), 
        .Q(\stage_3_retimer[6][16] ) );
  DFQD1 \stage_3_retimer_reg[6][15]  ( .D(\stage_3_output[6][15] ), .CP(clk), 
        .Q(\stage_3_retimer[6][15] ) );
  DFQD1 \stage_3_retimer_reg[6][14]  ( .D(\stage_3_output[6][14] ), .CP(clk), 
        .Q(\stage_3_retimer[6][14] ) );
  DFQD1 \stage_3_retimer_reg[6][13]  ( .D(\stage_3_output[6][13] ), .CP(clk), 
        .Q(\stage_3_retimer[6][13] ) );
  DFQD1 \stage_3_retimer_reg[6][12]  ( .D(\stage_3_output[6][12] ), .CP(clk), 
        .Q(\stage_3_retimer[6][12] ) );
  DFQD1 \stage_3_retimer_reg[6][11]  ( .D(\stage_3_output[6][11] ), .CP(clk), 
        .Q(\stage_3_retimer[6][11] ) );
  DFQD1 \stage_3_retimer_reg[6][10]  ( .D(\stage_3_output[6][10] ), .CP(clk), 
        .Q(\stage_3_retimer[6][10] ) );
  DFQD1 \stage_3_retimer_reg[6][9]  ( .D(\stage_3_output[6][9] ), .CP(clk), 
        .Q(\stage_3_retimer[6][9] ) );
  DFQD1 \stage_3_retimer_reg[6][8]  ( .D(\stage_3_output[6][8] ), .CP(clk), 
        .Q(\stage_3_retimer[6][8] ) );
  DFQD1 \stage_3_retimer_reg[6][7]  ( .D(\stage_3_output[6][7] ), .CP(clk), 
        .Q(\stage_3_retimer[6][7] ) );
  DFQD1 \stage_3_retimer_reg[6][6]  ( .D(\stage_3_output[6][6] ), .CP(clk), 
        .Q(\stage_3_retimer[6][6] ) );
  DFQD1 \stage_3_retimer_reg[6][5]  ( .D(\stage_3_output[6][5] ), .CP(clk), 
        .Q(\stage_3_retimer[6][5] ) );
  DFQD1 \stage_3_retimer_reg[6][4]  ( .D(\stage_3_output[6][4] ), .CP(clk), 
        .Q(\stage_3_retimer[6][4] ) );
  DFQD1 \stage_3_retimer_reg[6][3]  ( .D(\stage_3_output[6][3] ), .CP(clk), 
        .Q(\stage_3_retimer[6][3] ) );
  DFQD1 \stage_3_retimer_reg[6][2]  ( .D(\stage_3_output[6][2] ), .CP(clk), 
        .Q(\stage_3_retimer[6][2] ) );
  DFQD1 \stage_3_retimer_reg[6][1]  ( .D(\stage_3_output[6][1] ), .CP(clk), 
        .Q(\stage_3_retimer[6][1] ) );
  DFQD1 \stage_3_retimer_reg[6][0]  ( .D(\stage_3_output[6][0] ), .CP(clk), 
        .Q(\stage_3_retimer[6][0] ) );
  DFQD1 \stage_3_retimer_reg[5][19]  ( .D(\stage_3_output[5][19] ), .CP(clk), 
        .Q(\stage_3_retimer[5][19] ) );
  DFQD1 \stage_3_retimer_reg[5][18]  ( .D(\stage_3_output[5][18] ), .CP(clk), 
        .Q(\stage_3_retimer[5][18] ) );
  DFQD1 \stage_3_retimer_reg[5][17]  ( .D(\stage_3_output[5][17] ), .CP(clk), 
        .Q(\stage_3_retimer[5][17] ) );
  DFQD1 \stage_3_retimer_reg[5][16]  ( .D(\stage_3_output[5][16] ), .CP(clk), 
        .Q(\stage_3_retimer[5][16] ) );
  DFQD1 \stage_3_retimer_reg[5][15]  ( .D(\stage_3_output[5][15] ), .CP(clk), 
        .Q(\stage_3_retimer[5][15] ) );
  DFQD1 \stage_3_retimer_reg[5][14]  ( .D(\stage_3_output[5][14] ), .CP(clk), 
        .Q(\stage_3_retimer[5][14] ) );
  DFQD1 \stage_3_retimer_reg[5][13]  ( .D(\stage_3_output[5][13] ), .CP(clk), 
        .Q(\stage_3_retimer[5][13] ) );
  DFQD1 \stage_3_retimer_reg[5][12]  ( .D(\stage_3_output[5][12] ), .CP(clk), 
        .Q(\stage_3_retimer[5][12] ) );
  DFQD1 \stage_3_retimer_reg[5][11]  ( .D(\stage_3_output[5][11] ), .CP(clk), 
        .Q(\stage_3_retimer[5][11] ) );
  DFQD1 \stage_3_retimer_reg[5][10]  ( .D(\stage_3_output[5][10] ), .CP(clk), 
        .Q(\stage_3_retimer[5][10] ) );
  DFQD1 \stage_3_retimer_reg[5][9]  ( .D(\stage_3_output[5][9] ), .CP(clk), 
        .Q(\stage_3_retimer[5][9] ) );
  DFQD1 \stage_3_retimer_reg[5][8]  ( .D(\stage_3_output[5][8] ), .CP(clk), 
        .Q(\stage_3_retimer[5][8] ) );
  DFQD1 \stage_3_retimer_reg[5][7]  ( .D(\stage_3_output[5][7] ), .CP(clk), 
        .Q(\stage_3_retimer[5][7] ) );
  DFQD1 \stage_3_retimer_reg[5][6]  ( .D(\stage_3_output[5][6] ), .CP(clk), 
        .Q(\stage_3_retimer[5][6] ) );
  DFQD1 \stage_3_retimer_reg[5][5]  ( .D(\stage_3_output[5][5] ), .CP(clk), 
        .Q(\stage_3_retimer[5][5] ) );
  DFQD1 \stage_3_retimer_reg[5][4]  ( .D(\stage_3_output[5][4] ), .CP(clk), 
        .Q(\stage_3_retimer[5][4] ) );
  DFQD1 \stage_3_retimer_reg[5][3]  ( .D(\stage_3_output[5][3] ), .CP(clk), 
        .Q(\stage_3_retimer[5][3] ) );
  DFQD1 \stage_3_retimer_reg[5][2]  ( .D(\stage_3_output[5][2] ), .CP(clk), 
        .Q(\stage_3_retimer[5][2] ) );
  DFQD1 \stage_3_retimer_reg[5][1]  ( .D(\stage_3_output[5][1] ), .CP(clk), 
        .Q(\stage_3_retimer[5][1] ) );
  DFQD1 \stage_3_retimer_reg[5][0]  ( .D(\stage_3_output[5][0] ), .CP(clk), 
        .Q(\stage_3_retimer[5][0] ) );
  DFQD1 \stage_3_retimer_reg[4][19]  ( .D(\stage_3_output[4][19] ), .CP(clk), 
        .Q(\stage_3_retimer[4][19] ) );
  DFQD1 \stage_3_retimer_reg[4][18]  ( .D(\stage_3_output[4][18] ), .CP(clk), 
        .Q(\stage_3_retimer[4][18] ) );
  DFQD1 \stage_3_retimer_reg[4][17]  ( .D(\stage_3_output[4][17] ), .CP(clk), 
        .Q(\stage_3_retimer[4][17] ) );
  DFQD1 \stage_3_retimer_reg[4][16]  ( .D(\stage_3_output[4][16] ), .CP(clk), 
        .Q(\stage_3_retimer[4][16] ) );
  DFQD1 \stage_3_retimer_reg[4][15]  ( .D(\stage_3_output[4][15] ), .CP(clk), 
        .Q(\stage_3_retimer[4][15] ) );
  DFQD1 \stage_3_retimer_reg[4][14]  ( .D(\stage_3_output[4][14] ), .CP(clk), 
        .Q(\stage_3_retimer[4][14] ) );
  DFQD1 \stage_3_retimer_reg[4][13]  ( .D(\stage_3_output[4][13] ), .CP(clk), 
        .Q(\stage_3_retimer[4][13] ) );
  DFQD1 \stage_3_retimer_reg[4][12]  ( .D(\stage_3_output[4][12] ), .CP(clk), 
        .Q(\stage_3_retimer[4][12] ) );
  DFQD1 \stage_3_retimer_reg[4][11]  ( .D(\stage_3_output[4][11] ), .CP(clk), 
        .Q(\stage_3_retimer[4][11] ) );
  DFQD1 \stage_3_retimer_reg[4][10]  ( .D(\stage_3_output[4][10] ), .CP(clk), 
        .Q(\stage_3_retimer[4][10] ) );
  DFQD1 \stage_3_retimer_reg[4][9]  ( .D(\stage_3_output[4][9] ), .CP(clk), 
        .Q(\stage_3_retimer[4][9] ) );
  DFQD1 \stage_3_retimer_reg[4][8]  ( .D(\stage_3_output[4][8] ), .CP(clk), 
        .Q(\stage_3_retimer[4][8] ) );
  DFQD1 \stage_3_retimer_reg[4][7]  ( .D(\stage_3_output[4][7] ), .CP(clk), 
        .Q(\stage_3_retimer[4][7] ) );
  DFQD1 \stage_3_retimer_reg[4][6]  ( .D(\stage_3_output[4][6] ), .CP(clk), 
        .Q(\stage_3_retimer[4][6] ) );
  DFQD1 \stage_3_retimer_reg[4][5]  ( .D(\stage_3_output[4][5] ), .CP(clk), 
        .Q(\stage_3_retimer[4][5] ) );
  DFQD1 \stage_3_retimer_reg[4][4]  ( .D(\stage_3_output[4][4] ), .CP(clk), 
        .Q(\stage_3_retimer[4][4] ) );
  DFQD1 \stage_3_retimer_reg[4][3]  ( .D(\stage_3_output[4][3] ), .CP(clk), 
        .Q(\stage_3_retimer[4][3] ) );
  DFQD1 \stage_3_retimer_reg[4][2]  ( .D(\stage_3_output[4][2] ), .CP(clk), 
        .Q(\stage_3_retimer[4][2] ) );
  DFQD1 \stage_3_retimer_reg[4][1]  ( .D(\stage_3_output[4][1] ), .CP(clk), 
        .Q(\stage_3_retimer[4][1] ) );
  DFQD1 \stage_3_retimer_reg[4][0]  ( .D(\stage_3_output[4][0] ), .CP(clk), 
        .Q(\stage_3_retimer[4][0] ) );
  DFQD1 \stage_3_retimer_reg[3][19]  ( .D(\stage_3_output[3][19] ), .CP(clk), 
        .Q(\stage_3_retimer[3][19] ) );
  DFQD1 \stage_3_retimer_reg[3][18]  ( .D(\stage_3_output[3][18] ), .CP(clk), 
        .Q(\stage_3_retimer[3][18] ) );
  DFQD1 \stage_3_retimer_reg[3][17]  ( .D(\stage_3_output[3][17] ), .CP(clk), 
        .Q(\stage_3_retimer[3][17] ) );
  DFQD1 \stage_3_retimer_reg[3][16]  ( .D(\stage_3_output[3][16] ), .CP(clk), 
        .Q(\stage_3_retimer[3][16] ) );
  DFQD1 \stage_3_retimer_reg[3][15]  ( .D(\stage_3_output[3][15] ), .CP(clk), 
        .Q(\stage_3_retimer[3][15] ) );
  DFQD1 \stage_3_retimer_reg[3][14]  ( .D(\stage_3_output[3][14] ), .CP(clk), 
        .Q(\stage_3_retimer[3][14] ) );
  DFQD1 \stage_3_retimer_reg[3][13]  ( .D(\stage_3_output[3][13] ), .CP(clk), 
        .Q(\stage_3_retimer[3][13] ) );
  DFQD1 \stage_3_retimer_reg[3][12]  ( .D(\stage_3_output[3][12] ), .CP(clk), 
        .Q(\stage_3_retimer[3][12] ) );
  DFQD1 \stage_3_retimer_reg[3][11]  ( .D(\stage_3_output[3][11] ), .CP(clk), 
        .Q(\stage_3_retimer[3][11] ) );
  DFQD1 \stage_3_retimer_reg[3][10]  ( .D(\stage_3_output[3][10] ), .CP(clk), 
        .Q(\stage_3_retimer[3][10] ) );
  DFQD1 \stage_3_retimer_reg[3][9]  ( .D(\stage_3_output[3][9] ), .CP(clk), 
        .Q(\stage_3_retimer[3][9] ) );
  DFQD1 \stage_3_retimer_reg[3][8]  ( .D(\stage_3_output[3][8] ), .CP(clk), 
        .Q(\stage_3_retimer[3][8] ) );
  DFQD1 \stage_3_retimer_reg[3][7]  ( .D(\stage_3_output[3][7] ), .CP(clk), 
        .Q(\stage_3_retimer[3][7] ) );
  DFQD1 \stage_3_retimer_reg[3][6]  ( .D(\stage_3_output[3][6] ), .CP(clk), 
        .Q(\stage_3_retimer[3][6] ) );
  DFQD1 \stage_3_retimer_reg[3][5]  ( .D(\stage_3_output[3][5] ), .CP(clk), 
        .Q(\stage_3_retimer[3][5] ) );
  DFQD1 \stage_3_retimer_reg[3][4]  ( .D(\stage_3_output[3][4] ), .CP(clk), 
        .Q(\stage_3_retimer[3][4] ) );
  DFQD1 \stage_3_retimer_reg[3][3]  ( .D(\stage_3_output[3][3] ), .CP(clk), 
        .Q(\stage_3_retimer[3][3] ) );
  DFQD1 \stage_3_retimer_reg[3][2]  ( .D(\stage_3_output[3][2] ), .CP(clk), 
        .Q(\stage_3_retimer[3][2] ) );
  DFQD1 \stage_3_retimer_reg[3][1]  ( .D(\stage_3_output[3][1] ), .CP(clk), 
        .Q(\stage_3_retimer[3][1] ) );
  DFQD1 \stage_3_retimer_reg[3][0]  ( .D(\stage_3_output[3][0] ), .CP(clk), 
        .Q(\stage_3_retimer[3][0] ) );
  DFQD1 \stage_3_retimer_reg[2][19]  ( .D(\stage_3_output[2][19] ), .CP(clk), 
        .Q(\stage_3_retimer[2][19] ) );
  DFQD1 \stage_3_retimer_reg[2][18]  ( .D(\stage_3_output[2][18] ), .CP(clk), 
        .Q(\stage_3_retimer[2][18] ) );
  DFQD1 \stage_3_retimer_reg[2][17]  ( .D(\stage_3_output[2][17] ), .CP(clk), 
        .Q(\stage_3_retimer[2][17] ) );
  DFQD1 \stage_3_retimer_reg[2][16]  ( .D(\stage_3_output[2][16] ), .CP(clk), 
        .Q(\stage_3_retimer[2][16] ) );
  DFQD1 \stage_3_retimer_reg[2][15]  ( .D(\stage_3_output[2][15] ), .CP(clk), 
        .Q(\stage_3_retimer[2][15] ) );
  DFQD1 \stage_3_retimer_reg[2][14]  ( .D(\stage_3_output[2][14] ), .CP(clk), 
        .Q(\stage_3_retimer[2][14] ) );
  DFQD1 \stage_3_retimer_reg[2][13]  ( .D(\stage_3_output[2][13] ), .CP(clk), 
        .Q(\stage_3_retimer[2][13] ) );
  DFQD1 \stage_3_retimer_reg[2][12]  ( .D(\stage_3_output[2][12] ), .CP(clk), 
        .Q(\stage_3_retimer[2][12] ) );
  DFQD1 \stage_3_retimer_reg[2][11]  ( .D(\stage_3_output[2][11] ), .CP(clk), 
        .Q(\stage_3_retimer[2][11] ) );
  DFQD1 \stage_3_retimer_reg[2][10]  ( .D(\stage_3_output[2][10] ), .CP(clk), 
        .Q(\stage_3_retimer[2][10] ) );
  DFQD1 \stage_3_retimer_reg[2][9]  ( .D(\stage_3_output[2][9] ), .CP(clk), 
        .Q(\stage_3_retimer[2][9] ) );
  DFQD1 \stage_3_retimer_reg[2][8]  ( .D(\stage_3_output[2][8] ), .CP(clk), 
        .Q(\stage_3_retimer[2][8] ) );
  DFQD1 \stage_3_retimer_reg[2][7]  ( .D(\stage_3_output[2][7] ), .CP(clk), 
        .Q(\stage_3_retimer[2][7] ) );
  DFQD1 \stage_3_retimer_reg[2][6]  ( .D(\stage_3_output[2][6] ), .CP(clk), 
        .Q(\stage_3_retimer[2][6] ) );
  DFQD1 \stage_3_retimer_reg[2][5]  ( .D(\stage_3_output[2][5] ), .CP(clk), 
        .Q(\stage_3_retimer[2][5] ) );
  DFQD1 \stage_3_retimer_reg[2][4]  ( .D(\stage_3_output[2][4] ), .CP(clk), 
        .Q(\stage_3_retimer[2][4] ) );
  DFQD1 \stage_3_retimer_reg[2][3]  ( .D(\stage_3_output[2][3] ), .CP(clk), 
        .Q(\stage_3_retimer[2][3] ) );
  DFQD1 \stage_3_retimer_reg[2][2]  ( .D(\stage_3_output[2][2] ), .CP(clk), 
        .Q(\stage_3_retimer[2][2] ) );
  DFQD1 \stage_3_retimer_reg[2][1]  ( .D(\stage_3_output[2][1] ), .CP(clk), 
        .Q(\stage_3_retimer[2][1] ) );
  DFQD1 \stage_3_retimer_reg[2][0]  ( .D(\stage_3_output[2][0] ), .CP(clk), 
        .Q(\stage_3_retimer[2][0] ) );
  DFQD1 \stage_3_retimer_reg[1][19]  ( .D(\stage_3_output[1][19] ), .CP(clk), 
        .Q(\stage_3_retimer[1][19] ) );
  DFQD1 \stage_3_retimer_reg[1][18]  ( .D(\stage_3_output[1][18] ), .CP(clk), 
        .Q(\stage_3_retimer[1][18] ) );
  DFQD1 \stage_3_retimer_reg[1][17]  ( .D(\stage_3_output[1][17] ), .CP(clk), 
        .Q(\stage_3_retimer[1][17] ) );
  DFQD1 \stage_3_retimer_reg[1][16]  ( .D(\stage_3_output[1][16] ), .CP(clk), 
        .Q(\stage_3_retimer[1][16] ) );
  DFQD1 \stage_3_retimer_reg[1][15]  ( .D(\stage_3_output[1][15] ), .CP(clk), 
        .Q(\stage_3_retimer[1][15] ) );
  DFQD1 \stage_3_retimer_reg[1][14]  ( .D(\stage_3_output[1][14] ), .CP(clk), 
        .Q(\stage_3_retimer[1][14] ) );
  DFQD1 \stage_3_retimer_reg[1][13]  ( .D(\stage_3_output[1][13] ), .CP(clk), 
        .Q(\stage_3_retimer[1][13] ) );
  DFQD1 \stage_3_retimer_reg[1][12]  ( .D(\stage_3_output[1][12] ), .CP(clk), 
        .Q(\stage_3_retimer[1][12] ) );
  DFQD1 \stage_3_retimer_reg[1][11]  ( .D(\stage_3_output[1][11] ), .CP(clk), 
        .Q(\stage_3_retimer[1][11] ) );
  DFQD1 \stage_3_retimer_reg[1][10]  ( .D(\stage_3_output[1][10] ), .CP(clk), 
        .Q(\stage_3_retimer[1][10] ) );
  DFQD1 \stage_3_retimer_reg[1][9]  ( .D(\stage_3_output[1][9] ), .CP(clk), 
        .Q(\stage_3_retimer[1][9] ) );
  DFQD1 \stage_3_retimer_reg[1][8]  ( .D(\stage_3_output[1][8] ), .CP(clk), 
        .Q(\stage_3_retimer[1][8] ) );
  DFQD1 \stage_3_retimer_reg[1][7]  ( .D(\stage_3_output[1][7] ), .CP(clk), 
        .Q(\stage_3_retimer[1][7] ) );
  DFQD1 \stage_3_retimer_reg[1][6]  ( .D(\stage_3_output[1][6] ), .CP(clk), 
        .Q(\stage_3_retimer[1][6] ) );
  DFQD1 \stage_3_retimer_reg[1][5]  ( .D(\stage_3_output[1][5] ), .CP(clk), 
        .Q(\stage_3_retimer[1][5] ) );
  DFQD1 \stage_3_retimer_reg[1][4]  ( .D(\stage_3_output[1][4] ), .CP(clk), 
        .Q(\stage_3_retimer[1][4] ) );
  DFQD1 \stage_3_retimer_reg[1][3]  ( .D(\stage_3_output[1][3] ), .CP(clk), 
        .Q(\stage_3_retimer[1][3] ) );
  DFQD1 \stage_3_retimer_reg[1][2]  ( .D(\stage_3_output[1][2] ), .CP(clk), 
        .Q(\stage_3_retimer[1][2] ) );
  DFQD1 \stage_3_retimer_reg[1][1]  ( .D(\stage_3_output[1][1] ), .CP(clk), 
        .Q(\stage_3_retimer[1][1] ) );
  DFQD1 \stage_3_retimer_reg[1][0]  ( .D(\stage_3_output[1][0] ), .CP(clk), 
        .Q(\stage_3_retimer[1][0] ) );
  DFQD1 \stage_3_retimer_reg[0][19]  ( .D(\stage_3_output[0][19] ), .CP(clk), 
        .Q(\stage_3_retimer[0][19] ) );
  DFQD1 \stage_3_retimer_reg[0][18]  ( .D(\stage_3_output[0][18] ), .CP(clk), 
        .Q(\stage_3_retimer[0][18] ) );
  DFQD1 \stage_3_retimer_reg[0][17]  ( .D(\stage_3_output[0][17] ), .CP(clk), 
        .Q(\stage_3_retimer[0][17] ) );
  DFQD1 \stage_3_retimer_reg[0][16]  ( .D(\stage_3_output[0][16] ), .CP(clk), 
        .Q(\stage_3_retimer[0][16] ) );
  DFQD1 \stage_3_retimer_reg[0][15]  ( .D(\stage_3_output[0][15] ), .CP(clk), 
        .Q(\stage_3_retimer[0][15] ) );
  DFQD1 \stage_3_retimer_reg[0][14]  ( .D(\stage_3_output[0][14] ), .CP(clk), 
        .Q(\stage_3_retimer[0][14] ) );
  DFQD1 \stage_3_retimer_reg[0][13]  ( .D(\stage_3_output[0][13] ), .CP(clk), 
        .Q(\stage_3_retimer[0][13] ) );
  DFQD1 \stage_3_retimer_reg[0][12]  ( .D(\stage_3_output[0][12] ), .CP(clk), 
        .Q(\stage_3_retimer[0][12] ) );
  DFQD1 \stage_3_retimer_reg[0][11]  ( .D(\stage_3_output[0][11] ), .CP(clk), 
        .Q(\stage_3_retimer[0][11] ) );
  DFQD1 \stage_3_retimer_reg[0][10]  ( .D(\stage_3_output[0][10] ), .CP(clk), 
        .Q(\stage_3_retimer[0][10] ) );
  DFQD1 \stage_3_retimer_reg[0][9]  ( .D(\stage_3_output[0][9] ), .CP(clk), 
        .Q(\stage_3_retimer[0][9] ) );
  DFQD1 \stage_3_retimer_reg[0][8]  ( .D(\stage_3_output[0][8] ), .CP(clk), 
        .Q(\stage_3_retimer[0][8] ) );
  DFQD1 \stage_3_retimer_reg[0][7]  ( .D(\stage_3_output[0][7] ), .CP(clk), 
        .Q(\stage_3_retimer[0][7] ) );
  DFQD1 \stage_3_retimer_reg[0][6]  ( .D(\stage_3_output[0][6] ), .CP(clk), 
        .Q(\stage_3_retimer[0][6] ) );
  DFQD1 \stage_3_retimer_reg[0][5]  ( .D(\stage_3_output[0][5] ), .CP(clk), 
        .Q(\stage_3_retimer[0][5] ) );
  DFQD1 \stage_3_retimer_reg[0][4]  ( .D(\stage_3_output[0][4] ), .CP(clk), 
        .Q(\stage_3_retimer[0][4] ) );
  DFQD1 \stage_3_retimer_reg[0][3]  ( .D(\stage_3_output[0][3] ), .CP(clk), 
        .Q(\stage_3_retimer[0][3] ) );
  DFQD1 \stage_3_retimer_reg[0][2]  ( .D(\stage_3_output[0][2] ), .CP(clk), 
        .Q(\stage_3_retimer[0][2] ) );
  DFQD1 \stage_3_retimer_reg[0][1]  ( .D(\stage_3_output[0][1] ), .CP(clk), 
        .Q(\stage_3_retimer[0][1] ) );
  DFQD1 \stage_3_retimer_reg[0][0]  ( .D(\stage_3_output[0][0] ), .CP(clk), 
        .Q(\stage_3_retimer[0][0] ) );
  DFQD1 \stage_4_retimer_reg[7][19]  ( .D(\stage_4_output[7][19] ), .CP(clk), 
        .Q(out_output[19]) );
  DFQD1 \stage_4_retimer_reg[7][18]  ( .D(\stage_4_output[7][18] ), .CP(clk), 
        .Q(out_output[18]) );
  DFQD1 \stage_4_retimer_reg[7][17]  ( .D(\stage_4_output[7][17] ), .CP(clk), 
        .Q(out_output[17]) );
  DFQD1 \stage_4_retimer_reg[7][16]  ( .D(\stage_4_output[7][16] ), .CP(clk), 
        .Q(out_output[16]) );
  DFQD1 \stage_4_retimer_reg[7][15]  ( .D(\stage_4_output[7][15] ), .CP(clk), 
        .Q(out_output[15]) );
  DFQD1 \stage_4_retimer_reg[7][14]  ( .D(\stage_4_output[7][14] ), .CP(clk), 
        .Q(out_output[14]) );
  DFQD1 \stage_4_retimer_reg[7][13]  ( .D(\stage_4_output[7][13] ), .CP(clk), 
        .Q(out_output[13]) );
  DFQD1 \stage_4_retimer_reg[7][12]  ( .D(\stage_4_output[7][12] ), .CP(clk), 
        .Q(out_output[12]) );
  DFQD1 \stage_4_retimer_reg[7][11]  ( .D(\stage_4_output[7][11] ), .CP(clk), 
        .Q(out_output[11]) );
  DFQD1 \stage_4_retimer_reg[7][10]  ( .D(\stage_4_output[7][10] ), .CP(clk), 
        .Q(out_output[10]) );
  DFQD1 \stage_4_retimer_reg[7][9]  ( .D(\stage_4_output[7][9] ), .CP(clk), 
        .Q(out_output[9]) );
  DFQD1 \stage_4_retimer_reg[7][8]  ( .D(\stage_4_output[7][8] ), .CP(clk), 
        .Q(out_output[8]) );
  DFQD1 \stage_4_retimer_reg[7][7]  ( .D(\stage_4_output[7][7] ), .CP(clk), 
        .Q(out_output[7]) );
  DFQD1 \stage_4_retimer_reg[7][6]  ( .D(\stage_4_output[7][6] ), .CP(clk), 
        .Q(out_output[6]) );
  DFQD1 \stage_4_retimer_reg[7][5]  ( .D(\stage_4_output[7][5] ), .CP(clk), 
        .Q(out_output[5]) );
  DFQD1 \stage_4_retimer_reg[7][4]  ( .D(\stage_4_output[7][4] ), .CP(clk), 
        .Q(out_output[4]) );
  DFQD1 \stage_4_retimer_reg[7][3]  ( .D(\stage_4_output[7][3] ), .CP(clk), 
        .Q(out_output[3]) );
  DFQD1 \stage_4_retimer_reg[7][2]  ( .D(\stage_4_output[7][2] ), .CP(clk), 
        .Q(out_output[2]) );
  DFQD1 \stage_4_retimer_reg[7][1]  ( .D(\stage_4_output[7][1] ), .CP(clk), 
        .Q(out_output[1]) );
  DFQD1 \stage_4_retimer_reg[7][0]  ( .D(\stage_4_output[7][0] ), .CP(clk), 
        .Q(out_output[0]) );
  DFQD1 \stage_4_retimer_reg[6][19]  ( .D(\stage_4_output[6][19] ), .CP(clk), 
        .Q(out_output[39]) );
  DFQD1 \stage_4_retimer_reg[6][18]  ( .D(\stage_4_output[6][18] ), .CP(clk), 
        .Q(out_output[38]) );
  DFQD1 \stage_4_retimer_reg[6][17]  ( .D(\stage_4_output[6][17] ), .CP(clk), 
        .Q(out_output[37]) );
  DFQD1 \stage_4_retimer_reg[6][16]  ( .D(\stage_4_output[6][16] ), .CP(clk), 
        .Q(out_output[36]) );
  DFQD1 \stage_4_retimer_reg[6][15]  ( .D(\stage_4_output[6][15] ), .CP(clk), 
        .Q(out_output[35]) );
  DFQD1 \stage_4_retimer_reg[6][14]  ( .D(\stage_4_output[6][14] ), .CP(clk), 
        .Q(out_output[34]) );
  DFQD1 \stage_4_retimer_reg[6][13]  ( .D(\stage_4_output[6][13] ), .CP(clk), 
        .Q(out_output[33]) );
  DFQD1 \stage_4_retimer_reg[6][12]  ( .D(\stage_4_output[6][12] ), .CP(clk), 
        .Q(out_output[32]) );
  DFQD1 \stage_4_retimer_reg[6][11]  ( .D(\stage_4_output[6][11] ), .CP(clk), 
        .Q(out_output[31]) );
  DFQD1 \stage_4_retimer_reg[6][10]  ( .D(\stage_4_output[6][10] ), .CP(clk), 
        .Q(out_output[30]) );
  DFQD1 \stage_4_retimer_reg[6][9]  ( .D(\stage_4_output[6][9] ), .CP(clk), 
        .Q(out_output[29]) );
  DFQD1 \stage_4_retimer_reg[6][8]  ( .D(\stage_4_output[6][8] ), .CP(clk), 
        .Q(out_output[28]) );
  DFQD1 \stage_4_retimer_reg[6][7]  ( .D(\stage_4_output[6][7] ), .CP(clk), 
        .Q(out_output[27]) );
  DFQD1 \stage_4_retimer_reg[6][6]  ( .D(\stage_4_output[6][6] ), .CP(clk), 
        .Q(out_output[26]) );
  DFQD1 \stage_4_retimer_reg[6][5]  ( .D(\stage_4_output[6][5] ), .CP(clk), 
        .Q(out_output[25]) );
  DFQD1 \stage_4_retimer_reg[6][4]  ( .D(\stage_4_output[6][4] ), .CP(clk), 
        .Q(out_output[24]) );
  DFQD1 \stage_4_retimer_reg[6][3]  ( .D(\stage_4_output[6][3] ), .CP(clk), 
        .Q(out_output[23]) );
  DFQD1 \stage_4_retimer_reg[6][2]  ( .D(\stage_4_output[6][2] ), .CP(clk), 
        .Q(out_output[22]) );
  DFQD1 \stage_4_retimer_reg[6][1]  ( .D(\stage_4_output[6][1] ), .CP(clk), 
        .Q(out_output[21]) );
  DFQD1 \stage_4_retimer_reg[6][0]  ( .D(\stage_4_output[6][0] ), .CP(clk), 
        .Q(out_output[20]) );
  DFQD1 \stage_4_retimer_reg[5][19]  ( .D(\stage_4_output[5][19] ), .CP(clk), 
        .Q(out_output[59]) );
  DFQD1 \stage_4_retimer_reg[5][18]  ( .D(\stage_4_output[5][18] ), .CP(clk), 
        .Q(out_output[58]) );
  DFQD1 \stage_4_retimer_reg[5][17]  ( .D(\stage_4_output[5][17] ), .CP(clk), 
        .Q(out_output[57]) );
  DFQD1 \stage_4_retimer_reg[5][16]  ( .D(\stage_4_output[5][16] ), .CP(clk), 
        .Q(out_output[56]) );
  DFQD1 \stage_4_retimer_reg[5][15]  ( .D(\stage_4_output[5][15] ), .CP(clk), 
        .Q(out_output[55]) );
  DFQD1 \stage_4_retimer_reg[5][14]  ( .D(\stage_4_output[5][14] ), .CP(clk), 
        .Q(out_output[54]) );
  DFQD1 \stage_4_retimer_reg[5][13]  ( .D(\stage_4_output[5][13] ), .CP(clk), 
        .Q(out_output[53]) );
  DFQD1 \stage_4_retimer_reg[5][12]  ( .D(\stage_4_output[5][12] ), .CP(clk), 
        .Q(out_output[52]) );
  DFQD1 \stage_4_retimer_reg[5][11]  ( .D(\stage_4_output[5][11] ), .CP(clk), 
        .Q(out_output[51]) );
  DFQD1 \stage_4_retimer_reg[5][10]  ( .D(\stage_4_output[5][10] ), .CP(clk), 
        .Q(out_output[50]) );
  DFQD1 \stage_4_retimer_reg[5][9]  ( .D(\stage_4_output[5][9] ), .CP(clk), 
        .Q(out_output[49]) );
  DFQD1 \stage_4_retimer_reg[5][8]  ( .D(\stage_4_output[5][8] ), .CP(clk), 
        .Q(out_output[48]) );
  DFQD1 \stage_4_retimer_reg[5][7]  ( .D(\stage_4_output[5][7] ), .CP(clk), 
        .Q(out_output[47]) );
  DFQD1 \stage_4_retimer_reg[5][6]  ( .D(\stage_4_output[5][6] ), .CP(clk), 
        .Q(out_output[46]) );
  DFQD1 \stage_4_retimer_reg[5][5]  ( .D(\stage_4_output[5][5] ), .CP(clk), 
        .Q(out_output[45]) );
  DFQD1 \stage_4_retimer_reg[5][4]  ( .D(\stage_4_output[5][4] ), .CP(clk), 
        .Q(out_output[44]) );
  DFQD1 \stage_4_retimer_reg[5][3]  ( .D(\stage_4_output[5][3] ), .CP(clk), 
        .Q(out_output[43]) );
  DFQD1 \stage_4_retimer_reg[5][2]  ( .D(\stage_4_output[5][2] ), .CP(clk), 
        .Q(out_output[42]) );
  DFQD1 \stage_4_retimer_reg[5][1]  ( .D(\stage_4_output[5][1] ), .CP(clk), 
        .Q(out_output[41]) );
  DFQD1 \stage_4_retimer_reg[5][0]  ( .D(\stage_4_output[5][0] ), .CP(clk), 
        .Q(out_output[40]) );
  DFQD1 \stage_4_retimer_reg[4][19]  ( .D(\stage_4_output[4][19] ), .CP(clk), 
        .Q(out_output[79]) );
  DFQD1 \stage_4_retimer_reg[4][18]  ( .D(\stage_4_output[4][18] ), .CP(clk), 
        .Q(out_output[78]) );
  DFQD1 \stage_4_retimer_reg[4][17]  ( .D(\stage_4_output[4][17] ), .CP(clk), 
        .Q(out_output[77]) );
  DFQD1 \stage_4_retimer_reg[4][16]  ( .D(\stage_4_output[4][16] ), .CP(clk), 
        .Q(out_output[76]) );
  DFQD1 \stage_4_retimer_reg[4][15]  ( .D(\stage_4_output[4][15] ), .CP(clk), 
        .Q(out_output[75]) );
  DFQD1 \stage_4_retimer_reg[4][14]  ( .D(\stage_4_output[4][14] ), .CP(clk), 
        .Q(out_output[74]) );
  DFQD1 \stage_4_retimer_reg[4][13]  ( .D(\stage_4_output[4][13] ), .CP(clk), 
        .Q(out_output[73]) );
  DFQD1 \stage_4_retimer_reg[4][12]  ( .D(\stage_4_output[4][12] ), .CP(clk), 
        .Q(out_output[72]) );
  DFQD1 \stage_4_retimer_reg[4][11]  ( .D(\stage_4_output[4][11] ), .CP(clk), 
        .Q(out_output[71]) );
  DFQD1 \stage_4_retimer_reg[4][10]  ( .D(\stage_4_output[4][10] ), .CP(clk), 
        .Q(out_output[70]) );
  DFQD1 \stage_4_retimer_reg[4][9]  ( .D(\stage_4_output[4][9] ), .CP(clk), 
        .Q(out_output[69]) );
  DFQD1 \stage_4_retimer_reg[4][8]  ( .D(\stage_4_output[4][8] ), .CP(clk), 
        .Q(out_output[68]) );
  DFQD1 \stage_4_retimer_reg[4][7]  ( .D(\stage_4_output[4][7] ), .CP(clk), 
        .Q(out_output[67]) );
  DFQD1 \stage_4_retimer_reg[4][6]  ( .D(\stage_4_output[4][6] ), .CP(clk), 
        .Q(out_output[66]) );
  DFQD1 \stage_4_retimer_reg[4][5]  ( .D(\stage_4_output[4][5] ), .CP(clk), 
        .Q(out_output[65]) );
  DFQD1 \stage_4_retimer_reg[4][4]  ( .D(\stage_4_output[4][4] ), .CP(clk), 
        .Q(out_output[64]) );
  DFQD1 \stage_4_retimer_reg[4][3]  ( .D(\stage_4_output[4][3] ), .CP(clk), 
        .Q(out_output[63]) );
  DFQD1 \stage_4_retimer_reg[4][2]  ( .D(\stage_4_output[4][2] ), .CP(clk), 
        .Q(out_output[62]) );
  DFQD1 \stage_4_retimer_reg[4][1]  ( .D(\stage_4_output[4][1] ), .CP(clk), 
        .Q(out_output[61]) );
  DFQD1 \stage_4_retimer_reg[4][0]  ( .D(\stage_4_output[4][0] ), .CP(clk), 
        .Q(out_output[60]) );
  DFQD1 \stage_4_retimer_reg[3][19]  ( .D(\stage_4_output[3][19] ), .CP(clk), 
        .Q(out_output[99]) );
  DFQD1 \stage_4_retimer_reg[3][18]  ( .D(\stage_4_output[3][18] ), .CP(clk), 
        .Q(out_output[98]) );
  DFQD1 \stage_4_retimer_reg[3][17]  ( .D(\stage_4_output[3][17] ), .CP(clk), 
        .Q(out_output[97]) );
  DFQD1 \stage_4_retimer_reg[3][16]  ( .D(\stage_4_output[3][16] ), .CP(clk), 
        .Q(out_output[96]) );
  DFQD1 \stage_4_retimer_reg[3][15]  ( .D(\stage_4_output[3][15] ), .CP(clk), 
        .Q(out_output[95]) );
  DFQD1 \stage_4_retimer_reg[3][14]  ( .D(\stage_4_output[3][14] ), .CP(clk), 
        .Q(out_output[94]) );
  DFQD1 \stage_4_retimer_reg[3][13]  ( .D(\stage_4_output[3][13] ), .CP(clk), 
        .Q(out_output[93]) );
  DFQD1 \stage_4_retimer_reg[3][12]  ( .D(\stage_4_output[3][12] ), .CP(clk), 
        .Q(out_output[92]) );
  DFQD1 \stage_4_retimer_reg[3][11]  ( .D(\stage_4_output[3][11] ), .CP(clk), 
        .Q(out_output[91]) );
  DFQD1 \stage_4_retimer_reg[3][10]  ( .D(\stage_4_output[3][10] ), .CP(clk), 
        .Q(out_output[90]) );
  DFQD1 \stage_4_retimer_reg[3][9]  ( .D(\stage_4_output[3][9] ), .CP(clk), 
        .Q(out_output[89]) );
  DFQD1 \stage_4_retimer_reg[3][8]  ( .D(\stage_4_output[3][8] ), .CP(clk), 
        .Q(out_output[88]) );
  DFQD1 \stage_4_retimer_reg[3][7]  ( .D(\stage_4_output[3][7] ), .CP(clk), 
        .Q(out_output[87]) );
  DFQD1 \stage_4_retimer_reg[3][6]  ( .D(\stage_4_output[3][6] ), .CP(clk), 
        .Q(out_output[86]) );
  DFQD1 \stage_4_retimer_reg[3][5]  ( .D(\stage_4_output[3][5] ), .CP(clk), 
        .Q(out_output[85]) );
  DFQD1 \stage_4_retimer_reg[3][4]  ( .D(\stage_4_output[3][4] ), .CP(clk), 
        .Q(out_output[84]) );
  DFQD1 \stage_4_retimer_reg[3][3]  ( .D(\stage_4_output[3][3] ), .CP(clk), 
        .Q(out_output[83]) );
  DFQD1 \stage_4_retimer_reg[3][2]  ( .D(\stage_4_output[3][2] ), .CP(clk), 
        .Q(out_output[82]) );
  DFQD1 \stage_4_retimer_reg[3][1]  ( .D(\stage_4_output[3][1] ), .CP(clk), 
        .Q(out_output[81]) );
  DFQD1 \stage_4_retimer_reg[3][0]  ( .D(\stage_4_output[3][0] ), .CP(clk), 
        .Q(out_output[80]) );
  DFQD1 \stage_4_retimer_reg[2][19]  ( .D(\stage_4_output[2][19] ), .CP(clk), 
        .Q(out_output[119]) );
  DFQD1 \stage_4_retimer_reg[2][18]  ( .D(\stage_4_output[2][18] ), .CP(clk), 
        .Q(out_output[118]) );
  DFQD1 \stage_4_retimer_reg[2][17]  ( .D(\stage_4_output[2][17] ), .CP(clk), 
        .Q(out_output[117]) );
  DFQD1 \stage_4_retimer_reg[2][16]  ( .D(\stage_4_output[2][16] ), .CP(clk), 
        .Q(out_output[116]) );
  DFQD1 \stage_4_retimer_reg[2][15]  ( .D(\stage_4_output[2][15] ), .CP(clk), 
        .Q(out_output[115]) );
  DFQD1 \stage_4_retimer_reg[2][14]  ( .D(\stage_4_output[2][14] ), .CP(clk), 
        .Q(out_output[114]) );
  DFQD1 \stage_4_retimer_reg[2][13]  ( .D(\stage_4_output[2][13] ), .CP(clk), 
        .Q(out_output[113]) );
  DFQD1 \stage_4_retimer_reg[2][12]  ( .D(\stage_4_output[2][12] ), .CP(clk), 
        .Q(out_output[112]) );
  DFQD1 \stage_4_retimer_reg[2][11]  ( .D(\stage_4_output[2][11] ), .CP(clk), 
        .Q(out_output[111]) );
  DFQD1 \stage_4_retimer_reg[2][10]  ( .D(\stage_4_output[2][10] ), .CP(clk), 
        .Q(out_output[110]) );
  DFQD1 \stage_4_retimer_reg[2][9]  ( .D(\stage_4_output[2][9] ), .CP(clk), 
        .Q(out_output[109]) );
  DFQD1 \stage_4_retimer_reg[2][8]  ( .D(\stage_4_output[2][8] ), .CP(clk), 
        .Q(out_output[108]) );
  DFQD1 \stage_4_retimer_reg[2][7]  ( .D(\stage_4_output[2][7] ), .CP(clk), 
        .Q(out_output[107]) );
  DFQD1 \stage_4_retimer_reg[2][6]  ( .D(\stage_4_output[2][6] ), .CP(clk), 
        .Q(out_output[106]) );
  DFQD1 \stage_4_retimer_reg[2][5]  ( .D(\stage_4_output[2][5] ), .CP(clk), 
        .Q(out_output[105]) );
  DFQD1 \stage_4_retimer_reg[2][4]  ( .D(\stage_4_output[2][4] ), .CP(clk), 
        .Q(out_output[104]) );
  DFQD1 \stage_4_retimer_reg[2][3]  ( .D(\stage_4_output[2][3] ), .CP(clk), 
        .Q(out_output[103]) );
  DFQD1 \stage_4_retimer_reg[2][2]  ( .D(\stage_4_output[2][2] ), .CP(clk), 
        .Q(out_output[102]) );
  DFQD1 \stage_4_retimer_reg[2][1]  ( .D(\stage_4_output[2][1] ), .CP(clk), 
        .Q(out_output[101]) );
  DFQD1 \stage_4_retimer_reg[2][0]  ( .D(\stage_4_output[2][0] ), .CP(clk), 
        .Q(out_output[100]) );
  DFQD1 \stage_4_retimer_reg[1][19]  ( .D(\stage_4_output[1][19] ), .CP(clk), 
        .Q(out_output[139]) );
  DFQD1 \stage_4_retimer_reg[1][18]  ( .D(\stage_4_output[1][18] ), .CP(clk), 
        .Q(out_output[138]) );
  DFQD1 \stage_4_retimer_reg[1][17]  ( .D(\stage_4_output[1][17] ), .CP(clk), 
        .Q(out_output[137]) );
  DFQD1 \stage_4_retimer_reg[1][16]  ( .D(\stage_4_output[1][16] ), .CP(clk), 
        .Q(out_output[136]) );
  DFQD1 \stage_4_retimer_reg[1][15]  ( .D(\stage_4_output[1][15] ), .CP(clk), 
        .Q(out_output[135]) );
  DFQD1 \stage_4_retimer_reg[1][14]  ( .D(\stage_4_output[1][14] ), .CP(clk), 
        .Q(out_output[134]) );
  DFQD1 \stage_4_retimer_reg[1][13]  ( .D(\stage_4_output[1][13] ), .CP(clk), 
        .Q(out_output[133]) );
  DFQD1 \stage_4_retimer_reg[1][12]  ( .D(\stage_4_output[1][12] ), .CP(clk), 
        .Q(out_output[132]) );
  DFQD1 \stage_4_retimer_reg[1][11]  ( .D(\stage_4_output[1][11] ), .CP(clk), 
        .Q(out_output[131]) );
  DFQD1 \stage_4_retimer_reg[1][10]  ( .D(\stage_4_output[1][10] ), .CP(clk), 
        .Q(out_output[130]) );
  DFQD1 \stage_4_retimer_reg[1][9]  ( .D(\stage_4_output[1][9] ), .CP(clk), 
        .Q(out_output[129]) );
  DFQD1 \stage_4_retimer_reg[1][8]  ( .D(\stage_4_output[1][8] ), .CP(clk), 
        .Q(out_output[128]) );
  DFQD1 \stage_4_retimer_reg[1][7]  ( .D(\stage_4_output[1][7] ), .CP(clk), 
        .Q(out_output[127]) );
  DFQD1 \stage_4_retimer_reg[1][6]  ( .D(\stage_4_output[1][6] ), .CP(clk), 
        .Q(out_output[126]) );
  DFQD1 \stage_4_retimer_reg[1][5]  ( .D(\stage_4_output[1][5] ), .CP(clk), 
        .Q(out_output[125]) );
  DFQD1 \stage_4_retimer_reg[1][4]  ( .D(\stage_4_output[1][4] ), .CP(clk), 
        .Q(out_output[124]) );
  DFQD1 \stage_4_retimer_reg[1][3]  ( .D(\stage_4_output[1][3] ), .CP(clk), 
        .Q(out_output[123]) );
  DFQD1 \stage_4_retimer_reg[1][2]  ( .D(\stage_4_output[1][2] ), .CP(clk), 
        .Q(out_output[122]) );
  DFQD1 \stage_4_retimer_reg[1][1]  ( .D(\stage_4_output[1][1] ), .CP(clk), 
        .Q(out_output[121]) );
  DFQD1 \stage_4_retimer_reg[1][0]  ( .D(\stage_4_output[1][0] ), .CP(clk), 
        .Q(out_output[120]) );
  DFQD1 \stage_4_retimer_reg[0][19]  ( .D(\stage_4_output[0][19] ), .CP(clk), 
        .Q(out_output[159]) );
  DFQD1 \stage_4_retimer_reg[0][18]  ( .D(\stage_4_output[0][18] ), .CP(clk), 
        .Q(out_output[158]) );
  DFQD1 \stage_4_retimer_reg[0][17]  ( .D(\stage_4_output[0][17] ), .CP(clk), 
        .Q(out_output[157]) );
  DFQD1 \stage_4_retimer_reg[0][16]  ( .D(\stage_4_output[0][16] ), .CP(clk), 
        .Q(out_output[156]) );
  DFQD1 \stage_4_retimer_reg[0][15]  ( .D(\stage_4_output[0][15] ), .CP(clk), 
        .Q(out_output[155]) );
  DFQD1 \stage_4_retimer_reg[0][14]  ( .D(\stage_4_output[0][14] ), .CP(clk), 
        .Q(out_output[154]) );
  DFQD1 \stage_4_retimer_reg[0][13]  ( .D(\stage_4_output[0][13] ), .CP(clk), 
        .Q(out_output[153]) );
  DFQD1 \stage_4_retimer_reg[0][12]  ( .D(\stage_4_output[0][12] ), .CP(clk), 
        .Q(out_output[152]) );
  DFQD1 \stage_4_retimer_reg[0][11]  ( .D(\stage_4_output[0][11] ), .CP(clk), 
        .Q(out_output[151]) );
  DFQD1 \stage_4_retimer_reg[0][10]  ( .D(\stage_4_output[0][10] ), .CP(clk), 
        .Q(out_output[150]) );
  DFQD1 \stage_4_retimer_reg[0][9]  ( .D(\stage_4_output[0][9] ), .CP(clk), 
        .Q(out_output[149]) );
  DFQD1 \stage_4_retimer_reg[0][8]  ( .D(\stage_4_output[0][8] ), .CP(clk), 
        .Q(out_output[148]) );
  DFQD1 \stage_4_retimer_reg[0][7]  ( .D(\stage_4_output[0][7] ), .CP(clk), 
        .Q(out_output[147]) );
  DFQD1 \stage_4_retimer_reg[0][6]  ( .D(\stage_4_output[0][6] ), .CP(clk), 
        .Q(out_output[146]) );
  DFQD1 \stage_4_retimer_reg[0][5]  ( .D(\stage_4_output[0][5] ), .CP(clk), 
        .Q(out_output[145]) );
  DFQD1 \stage_4_retimer_reg[0][4]  ( .D(\stage_4_output[0][4] ), .CP(clk), 
        .Q(out_output[144]) );
  DFQD1 \stage_4_retimer_reg[0][3]  ( .D(\stage_4_output[0][3] ), .CP(clk), 
        .Q(out_output[143]) );
  DFQD1 \stage_4_retimer_reg[0][2]  ( .D(\stage_4_output[0][2] ), .CP(clk), 
        .Q(out_output[142]) );
  DFQD1 \stage_4_retimer_reg[0][1]  ( .D(\stage_4_output[0][1] ), .CP(clk), 
        .Q(out_output[141]) );
  DFQD1 \stage_4_retimer_reg[0][0]  ( .D(\stage_4_output[0][0] ), .CP(clk), 
        .Q(out_output[140]) );
  TIEH U3 ( .Z(\*Logic1* ) );
endmodule

