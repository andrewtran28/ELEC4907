
module routing_engine ( port_dest, control, done, clk, rst );
  input [31:0] port_dest;
  output [19:0] control;
  input clk, rst;
  output done;
  wire   \dst[0][2] , \dst[0][1] , \dst[0][0] , \dst[1][2] , \dst[1][1] ,
         \dst[2][2] , \dst[2][1] , \dst[2][0] , \dst[3][2] , \dst[3][0] ,
         \dst[4][2] , \dst[4][1] , \dst[4][0] , \dst[5][2] , \dst[5][1] ,
         \dst[5][0] , \dst[6][2] , \dst[6][1] , \dst[6][0] , \dst[7][1] ,
         \dst[7][0] , N696, N697, N698, N699, N812, N813, N925, N926, N927,
         N1024, N1025, N1136, N1137, N1138, N1139, N1250, N1251, N1252, N1253,
         N1365, N1366, N1448, N1449, N1450, N1566, N1569, N1570, N1576, N1577,
         N1578, \stage_1_output[0][1] , \stage_1_output[0][2] ,
         \stage_1_output[1][2] , \stage_1_output[2][1] ,
         \stage_1_output[2][2] , \stage_1_output[3][2] ,
         \stage_1_output[4][1] , \stage_1_output[6][1] , N1614, N1615, N1616,
         N1618, n6, n865, n870, n1281, n1669, n1670, n1674, n1675, n1685,
         n1698, n1704, \control[13] , n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461;
  assign control[19] = \control[13] ;
  assign control[15] = \control[13] ;
  assign control[13] = \control[13] ;

  EDFQD1 \dst_reg[0][0]  ( .D(N697), .E(N696), .CP(clk), .Q(\dst[0][0] ) );
  EDFQD1 \dst_reg[1][2]  ( .D(N813), .E(n1704), .CP(clk), .Q(\dst[1][2] ) );
  EDFQD1 \dst_reg[1][1]  ( .D(N812), .E(n1704), .CP(clk), .Q(\dst[1][1] ) );
  EDFQD1 \dst_reg[5][2]  ( .D(N1253), .E(N1250), .CP(clk), .Q(\dst[5][2] ) );
  EDFQD1 \dst_reg[0][1]  ( .D(N698), .E(N696), .CP(clk), .Q(\dst[0][1] ) );
  EDFQD1 \dst_reg[0][2]  ( .D(N699), .E(N696), .CP(clk), .Q(\dst[0][2] ) );
  EDFQD1 \dst_reg[2][2]  ( .D(N927), .E(n1698), .CP(clk), .Q(\dst[2][2] ) );
  EDFQD1 \dst_reg[2][1]  ( .D(N926), .E(n1698), .CP(clk), .Q(\dst[2][1] ) );
  EDFQD1 \dst_reg[2][0]  ( .D(N925), .E(n1698), .CP(clk), .Q(\dst[2][0] ) );
  EDFQD1 \dst_reg[3][2]  ( .D(N1025), .E(n870), .CP(clk), .Q(\dst[3][2] ) );
  EDFQD1 \dst_reg[3][0]  ( .D(N1024), .E(n870), .CP(clk), .Q(\dst[3][0] ) );
  EDFQD1 \dst_reg[4][2]  ( .D(N1139), .E(N1136), .CP(clk), .Q(\dst[4][2] ) );
  EDFQD1 \dst_reg[4][1]  ( .D(N1138), .E(N1136), .CP(clk), .Q(\dst[4][1] ) );
  EDFQD1 \dst_reg[4][0]  ( .D(N1137), .E(N1136), .CP(clk), .Q(\dst[4][0] ) );
  EDFQD1 \dst_reg[5][1]  ( .D(N1252), .E(N1250), .CP(clk), .Q(\dst[5][1] ) );
  EDFQD1 \dst_reg[5][0]  ( .D(N1251), .E(N1250), .CP(clk), .Q(\dst[5][0] ) );
  EDFQD1 \dst_reg[7][1]  ( .D(N1450), .E(N1448), .CP(clk), .Q(\dst[7][1] ) );
  EDFQD1 \dst_reg[7][0]  ( .D(N1449), .E(N1448), .CP(clk), .Q(\dst[7][0] ) );
  EDFQD1 \dst_reg[6][1]  ( .D(N1366), .E(n2079), .CP(clk), .Q(\dst[6][1] ) );
  EDFQD1 \dst_reg[6][0]  ( .D(N1365), .E(n2079), .CP(clk), .Q(\dst[6][0] ) );
  EDFQD1 \dst_reg[6][2]  ( .D(n1685), .E(n2079), .CP(clk), .Q(\dst[6][2] ) );
  DFQD1 \stage_1_output_reg[4][1]  ( .D(N1569), .CP(clk), .Q(
        \stage_1_output[4][1] ) );
  DFQD1 \stage_1_output_reg[6][1]  ( .D(N1618), .CP(clk), .Q(
        \stage_1_output[6][1] ) );
  DFQD1 \stage_1_output_reg[0][1]  ( .D(n1675), .CP(clk), .Q(
        \stage_1_output[0][1] ) );
  DFQD1 \stage_1_output_reg[2][1]  ( .D(N1615), .CP(clk), .Q(
        \stage_1_output[2][1] ) );
  DFQD1 \stage_1_output_reg[0][2]  ( .D(N1566), .CP(clk), .Q(
        \stage_1_output[0][2] ) );
  DFQD1 \stage_1_output_reg[1][2]  ( .D(N1576), .CP(clk), .Q(
        \stage_1_output[1][2] ) );
  DFQD1 \stage_1_output_reg[2][2]  ( .D(N1614), .CP(clk), .Q(
        \stage_1_output[2][2] ) );
  DFQD1 \stage_1_output_reg[3][2]  ( .D(N1616), .CP(clk), .Q(
        \stage_1_output[3][2] ) );
  DFQD2 \stage_1_output_reg[4][0]  ( .D(N1570), .CP(clk), .Q(control[9]) );
  DFQD2 \stage_1_output_reg[1][0]  ( .D(N1577), .CP(clk), .Q(control[10]) );
  DFQD2 \stage_1_output_reg[0][0]  ( .D(n1674), .CP(clk), .Q(control[11]) );
  DFQD2 \stage_0_sw_ctl_reg[3]  ( .D(n6), .CP(clk), .Q(control[16]) );
  DFQD2 \stage_1_output_reg[5][0]  ( .D(N1578), .CP(clk), .Q(control[8]) );
  DFQD2 \stage_1_sw_ctl_reg[1]  ( .D(n1281), .CP(clk), .Q(control[14]) );
  DFQD2 \stage_1_sw_ctl_reg[3]  ( .D(n1670), .CP(clk), .Q(control[12]) );
  DFQD2 \stage_0_sw_ctl_reg[2]  ( .D(n865), .CP(clk), .Q(control[17]) );
  DFQD2 \stage_0_sw_ctl_reg[1]  ( .D(n1669), .CP(clk), .Q(control[18]) );
  MUX2ND2 U1426 ( .I0(n2083), .I1(n2084), .S(control[7]), .ZN(control[3]) );
  MUX2ND2 U1427 ( .I0(n2081), .I1(n2082), .S(control[9]), .ZN(control[5]) );
  MUX2ND2 U1428 ( .I0(n2084), .I1(n2083), .S(control[7]), .ZN(control[2]) );
  CKMUX2D2 U1429 ( .I0(\stage_1_output[0][1] ), .I1(\stage_1_output[2][1] ), 
        .S(control[11]), .Z(control[7]) );
  MUX2ND2 U1430 ( .I0(n2082), .I1(n2081), .S(control[9]), .ZN(control[4]) );
  MUX2ND2 U1431 ( .I0(n2086), .I1(n2085), .S(control[6]), .ZN(control[0]) );
  MUX2ND2 U1432 ( .I0(n2085), .I1(n2086), .S(control[6]), .ZN(control[1]) );
  CKMUX2D2 U1433 ( .I0(\stage_1_output[2][1] ), .I1(\stage_1_output[0][1] ), 
        .S(control[11]), .Z(control[6]) );
  TIEH U1434 ( .Z(done) );
  TIEL U1435 ( .ZN(\control[13] ) );
  CKND0 U1436 ( .I(n2080), .ZN(n2079) );
  CKND0 U1437 ( .I(\stage_1_output[4][1] ), .ZN(n2081) );
  CKND0 U1438 ( .I(\stage_1_output[6][1] ), .ZN(n2082) );
  MUX2ND0 U1439 ( .I0(\stage_1_output[0][2] ), .I1(\stage_1_output[2][2] ), 
        .S(control[11]), .ZN(n2083) );
  MUX2ND0 U1440 ( .I0(\stage_1_output[1][2] ), .I1(\stage_1_output[3][2] ), 
        .S(control[10]), .ZN(n2084) );
  MUX2ND0 U1441 ( .I0(\stage_1_output[2][2] ), .I1(\stage_1_output[0][2] ), 
        .S(control[11]), .ZN(n2085) );
  MUX2ND0 U1442 ( .I0(\stage_1_output[3][2] ), .I1(\stage_1_output[1][2] ), 
        .S(control[10]), .ZN(n2086) );
  MUX3ND0 U1443 ( .I0(n2087), .I1(n2088), .I2(n2089), .S0(n865), .S1(n1670), 
        .ZN(N1618) );
  CKXOR2D0 U1444 ( .A1(n2090), .A2(N1570), .Z(n1670) );
  MUX2ND0 U1445 ( .I0(n2091), .I1(n2092), .S(n865), .ZN(n2090) );
  MUX2D0 U1446 ( .I0(n2093), .I1(n2094), .S(n6), .Z(n2089) );
  MUX2ND0 U1447 ( .I0(n2095), .I1(n2096), .S(n2097), .ZN(N1616) );
  MUX3ND0 U1448 ( .I0(n2094), .I1(n2093), .I2(n2098), .S0(n6), .S1(n2097), 
        .ZN(N1615) );
  MUX2D0 U1449 ( .I0(n2088), .I1(n2087), .S(n865), .Z(n2098) );
  MUX2ND0 U1450 ( .I0(\dst[5][1] ), .I1(N1252), .S(N1250), .ZN(n2087) );
  MUX2ND0 U1451 ( .I0(\dst[7][1] ), .I1(N1450), .S(N1448), .ZN(n2093) );
  MUX2ND0 U1452 ( .I0(n2096), .I1(n2095), .S(n2097), .ZN(N1614) );
  CKND0 U1453 ( .I(n1281), .ZN(n2097) );
  CKXOR2D0 U1454 ( .A1(n2099), .A2(n1674), .Z(n1281) );
  MUX2ND0 U1455 ( .I0(n2092), .I1(n2091), .S(n865), .ZN(n2099) );
  MUX2D0 U1456 ( .I0(\dst[5][2] ), .I1(N1253), .S(N1250), .Z(n2091) );
  MUX2D0 U1457 ( .I0(n2100), .I1(n2101), .S(n865), .Z(n2095) );
  AN4D0 U1458 ( .A1(n2102), .A2(n2103), .A3(n2104), .A4(n2105), .Z(n865) );
  MUX2ND0 U1459 ( .I0(\dst[5][0] ), .I1(N1251), .S(N1250), .ZN(n2101) );
  MUX2ND0 U1460 ( .I0(\dst[4][0] ), .I1(N1137), .S(N1136), .ZN(n2100) );
  MUX2D0 U1461 ( .I0(n2106), .I1(n2107), .S(n6), .Z(n2096) );
  MUX3D0 U1462 ( .I0(n2108), .I1(n2109), .I2(n2110), .S0(n1685), .S1(n2080), 
        .Z(n6) );
  AO211D0 U1463 ( .A1(n2111), .A2(n2112), .B(n2113), .C(n2114), .Z(n1685) );
  AO21D0 U1464 ( .A1(n2115), .A2(port_dest[6]), .B(n2116), .Z(n2111) );
  MUX2D0 U1465 ( .I0(n2108), .I1(n2109), .S(\dst[6][2] ), .Z(n2110) );
  OAI21D0 U1466 ( .A1(n2117), .A2(n2118), .B(n2119), .ZN(n2109) );
  MUX2ND0 U1467 ( .I0(n2120), .I1(n2121), .S(n2094), .ZN(n2119) );
  CKND2D0 U1468 ( .A1(n2122), .A2(n2102), .ZN(n2121) );
  ND4D0 U1469 ( .A1(n2092), .A2(n2088), .A3(n2122), .A4(n2123), .ZN(n2102) );
  CKND2D0 U1470 ( .A1(n2124), .A2(n2103), .ZN(n2120) );
  ND4D0 U1471 ( .A1(n2125), .A2(n2092), .A3(n2124), .A4(n2126), .ZN(n2103) );
  CKND0 U1472 ( .I(n2127), .ZN(n2092) );
  OAI21D0 U1473 ( .A1(n1674), .A2(n2118), .B(n2128), .ZN(n2108) );
  MUX2ND0 U1474 ( .I0(n2129), .I1(n2130), .S(n2094), .ZN(n2128) );
  CKND2D0 U1475 ( .A1(n2131), .A2(n2104), .ZN(n2130) );
  ND4D0 U1476 ( .A1(n2127), .A2(n2088), .A3(n2131), .A4(n2132), .ZN(n2104) );
  CKND2D0 U1477 ( .A1(n2133), .A2(n2105), .ZN(n2129) );
  ND4D0 U1478 ( .A1(n2125), .A2(n2127), .A3(n2133), .A4(n2134), .ZN(n2105) );
  MUX2ND0 U1479 ( .I0(\dst[4][2] ), .I1(N1139), .S(N1136), .ZN(n2127) );
  CKND0 U1480 ( .I(n2088), .ZN(n2125) );
  MUX2ND0 U1481 ( .I0(\dst[4][1] ), .I1(N1138), .S(N1136), .ZN(n2088) );
  CKXOR2D0 U1482 ( .A1(n2094), .A2(n2135), .Z(n2118) );
  MUX2ND0 U1483 ( .I0(N1366), .I1(\dst[6][1] ), .S(n2080), .ZN(n2094) );
  MUX2ND0 U1484 ( .I0(\dst[7][0] ), .I1(N1449), .S(N1448), .ZN(n2107) );
  MUX2ND0 U1485 ( .I0(N1365), .I1(\dst[6][0] ), .S(n2080), .ZN(n2106) );
  IINR4D0 U1486 ( .A1(n2136), .A2(n2137), .B1(n2116), .B2(n2138), .ZN(n2080)
         );
  ND3D0 U1487 ( .A1(n2139), .A2(n2140), .A3(n2141), .ZN(n2116) );
  INR2D0 U1488 ( .A1(n2142), .B1(n2143), .ZN(n2136) );
  MUX2ND0 U1489 ( .I0(n2144), .I1(n2145), .S(n1669), .ZN(N1578) );
  MUX2ND0 U1490 ( .I0(n2145), .I1(n2144), .S(n1669), .ZN(N1577) );
  MUX2ND0 U1491 ( .I0(\dst[3][2] ), .I1(N1025), .S(n870), .ZN(n2144) );
  MUX2ND0 U1492 ( .I0(n2146), .I1(n2147), .S(n1669), .ZN(N1576) );
  AN4D0 U1493 ( .A1(n2122), .A2(n2124), .A3(n2131), .A4(n2133), .Z(n1669) );
  ND3D0 U1494 ( .A1(n2145), .A2(n2134), .A3(n2148), .ZN(n2133) );
  CKND2D0 U1495 ( .A1(n1675), .A2(n2117), .ZN(n2134) );
  ND3D0 U1496 ( .A1(n2145), .A2(n2132), .A3(n2149), .ZN(n2131) );
  CKND2D0 U1497 ( .A1(n2135), .A2(n2117), .ZN(n2132) );
  ND3D0 U1498 ( .A1(n2148), .A2(n2126), .A3(n2150), .ZN(n2124) );
  CKND2D0 U1499 ( .A1(n1674), .A2(n1675), .ZN(n2126) );
  CKND0 U1500 ( .I(n2135), .ZN(n1675) );
  CKND0 U1501 ( .I(n2149), .ZN(n2148) );
  ND3D0 U1502 ( .A1(n2149), .A2(n2123), .A3(n2150), .ZN(n2122) );
  CKND0 U1503 ( .I(n2145), .ZN(n2150) );
  MUX2ND0 U1504 ( .I0(\dst[2][2] ), .I1(N927), .S(n1698), .ZN(n2145) );
  OAI211D0 U1505 ( .A1(port_dest[23]), .A2(n2151), .B(n2152), .C(n2153), .ZN(
        N927) );
  AOI21D0 U1506 ( .A1(n2154), .A2(port_dest[22]), .B(n2155), .ZN(n2151) );
  CKND2D0 U1507 ( .A1(n1674), .A2(n2135), .ZN(n2123) );
  MUX2ND0 U1508 ( .I0(\dst[0][1] ), .I1(N698), .S(N696), .ZN(n2135) );
  OAI211D0 U1509 ( .A1(n2156), .A2(n2157), .B(n2158), .C(n2159), .ZN(N698) );
  MUX2ND0 U1510 ( .I0(n2160), .I1(port_dest[29]), .S(port_dest[31]), .ZN(n2159) );
  CKND2D0 U1511 ( .A1(n2161), .A2(n2162), .ZN(n2157) );
  AOI22D0 U1512 ( .A1(n2163), .A2(n2164), .B1(n2165), .B2(n2166), .ZN(n2156)
         );
  OAI21D0 U1513 ( .A1(port_dest[31]), .A2(n2167), .B(n2168), .ZN(n2164) );
  CKND0 U1514 ( .I(n2117), .ZN(n1674) );
  MUX2ND0 U1515 ( .I0(\dst[0][2] ), .I1(N699), .S(N696), .ZN(n2117) );
  OAI221D0 U1516 ( .A1(port_dest[31]), .A2(n2169), .B1(n2170), .B2(n2171), .C(
        n2172), .ZN(N699) );
  NR2D0 U1517 ( .A1(n2173), .A2(n2174), .ZN(n2172) );
  MUX2ND0 U1518 ( .I0(\dst[2][1] ), .I1(N926), .S(n1698), .ZN(n2149) );
  OAI221D0 U1519 ( .A1(n2175), .A2(n2176), .B1(port_dest[23]), .B2(n2177), .C(
        n2153), .ZN(N926) );
  INR2D0 U1520 ( .A1(n2178), .B1(n2179), .ZN(n2177) );
  AOI21D0 U1521 ( .A1(n2180), .A2(n2181), .B(port_dest[23]), .ZN(n2175) );
  MUX2ND0 U1522 ( .I0(\dst[3][0] ), .I1(N1024), .S(n870), .ZN(n2147) );
  IND2D0 U1523 ( .A1(n2182), .B1(n2183), .ZN(n870) );
  MUX2ND0 U1524 ( .I0(\dst[2][0] ), .I1(N925), .S(n1698), .ZN(n2146) );
  IND4D0 U1525 ( .A1(n2155), .B1(n2178), .B2(n2184), .B3(n2181), .ZN(n1698) );
  NR2D0 U1526 ( .A1(port_dest[23]), .A2(n2185), .ZN(n2184) );
  IAO21D0 U1527 ( .A1(n2186), .A2(n2187), .B(n2188), .ZN(n2178) );
  IND2D0 U1528 ( .A1(n2179), .B1(n2180), .ZN(n2155) );
  AOI22D0 U1529 ( .A1(n2154), .A2(n2189), .B1(n2190), .B2(n2191), .ZN(n2180)
         );
  CKND2D0 U1530 ( .A1(n2192), .A2(n2153), .ZN(N925) );
  IND2D0 U1531 ( .A1(n2193), .B1(n2185), .ZN(n2153) );
  MUX2ND0 U1532 ( .I0(n2194), .I1(port_dest[20]), .S(port_dest[23]), .ZN(n2192) );
  NR2D0 U1533 ( .A1(n2179), .A2(n2195), .ZN(n2194) );
  AOI22D0 U1534 ( .A1(n2196), .A2(n2197), .B1(n2191), .B2(n2190), .ZN(n2195)
         );
  CKND0 U1535 ( .I(n2198), .ZN(n2190) );
  OAI32D0 U1536 ( .A1(n2199), .A2(n2200), .A3(n2188), .B1(n2186), .B2(n2187), 
        .ZN(n2197) );
  INR2D0 U1537 ( .A1(n2181), .B1(n2201), .ZN(n2188) );
  NR2D0 U1538 ( .A1(n2202), .A2(port_dest[20]), .ZN(n2199) );
  CKND2D0 U1539 ( .A1(n2189), .A2(n2154), .ZN(n2196) );
  CKND0 U1540 ( .I(n2203), .ZN(n2189) );
  NR3D0 U1541 ( .A1(n2198), .A2(n2191), .A3(n2204), .ZN(n2179) );
  MUX2D0 U1542 ( .I0(\dst[1][2] ), .I1(N813), .S(n1704), .Z(N1570) );
  OAI211D0 U1543 ( .A1(n2205), .A2(n2206), .B(n2207), .C(n2208), .ZN(N813) );
  IAO21D0 U1544 ( .A1(n2209), .A2(port_dest[27]), .B(n2210), .ZN(n2208) );
  MUX2D0 U1545 ( .I0(\dst[1][1] ), .I1(N812), .S(n1704), .Z(N1569) );
  ND4D0 U1546 ( .A1(n2211), .A2(n2212), .A3(n2209), .A4(n2213), .ZN(n1704) );
  OAI221D0 U1547 ( .A1(n2214), .A2(n2215), .B1(n2216), .B2(n2217), .C(n2207), 
        .ZN(N812) );
  OA22D0 U1548 ( .A1(port_dest[27]), .A2(n2212), .B1(n2218), .B2(n2213), .Z(
        n2207) );
  ND4D0 U1549 ( .A1(n2219), .A2(n2220), .A3(n2221), .A4(n2222), .ZN(n2212) );
  AN2D0 U1550 ( .A1(n2216), .A2(n2223), .Z(n2222) );
  AOI21D0 U1551 ( .A1(n2221), .A2(n2209), .B(port_dest[27]), .ZN(n2214) );
  OAI211D0 U1552 ( .A1(n2224), .A2(n2225), .B(n2221), .C(n2216), .ZN(n2209) );
  MUX2D0 U1553 ( .I0(\dst[0][0] ), .I1(N697), .S(N696), .Z(N1566) );
  IND3D0 U1554 ( .A1(n2171), .B1(n2226), .B2(n2169), .ZN(N696) );
  AN3D0 U1555 ( .A1(n2227), .A2(n2161), .A3(n2162), .Z(n2169) );
  CKND2D0 U1556 ( .A1(n2228), .A2(n2158), .ZN(N697) );
  CKND0 U1557 ( .I(n2174), .ZN(n2158) );
  NR2D0 U1558 ( .A1(n2229), .A2(n2226), .ZN(n2174) );
  MUX2ND0 U1559 ( .I0(n2230), .I1(port_dest[28]), .S(port_dest[31]), .ZN(n2228) );
  AOI21D0 U1560 ( .A1(n2162), .A2(n2231), .B(n2160), .ZN(n2230) );
  CKND0 U1561 ( .I(n2227), .ZN(n2160) );
  IND4D0 U1562 ( .A1(n2232), .B1(n2233), .B2(n2234), .B3(n2235), .ZN(n2227) );
  NR2D0 U1563 ( .A1(n2166), .A2(n2236), .ZN(n2233) );
  CKND0 U1564 ( .I(n2237), .ZN(n2166) );
  CKND2D0 U1565 ( .A1(n2238), .A2(n2161), .ZN(n2231) );
  ND3D0 U1566 ( .A1(n2234), .A2(n2237), .A3(n2239), .ZN(n2161) );
  OAI22D0 U1567 ( .A1(n2240), .A2(n2237), .B1(n2241), .B2(n2242), .ZN(n2238)
         );
  AOI21D0 U1568 ( .A1(port_dest[28]), .A2(n2167), .B(n2243), .ZN(n2242) );
  ND4D0 U1569 ( .A1(n2236), .A2(n2234), .A3(n2235), .A4(n2237), .ZN(n2162) );
  CKND0 U1570 ( .I(n2240), .ZN(n2234) );
  CKND0 U1571 ( .I(n2244), .ZN(n2236) );
  CKND2D0 U1572 ( .A1(n2245), .A2(n2246), .ZN(N1450) );
  OAI31D0 U1573 ( .A1(n2247), .A2(n2248), .A3(n2249), .B(n2250), .ZN(n2246) );
  CKND0 U1574 ( .I(n2251), .ZN(n2248) );
  AOI211D0 U1575 ( .A1(n2252), .A2(n2253), .B(n2254), .C(n2255), .ZN(n2247) );
  CKND2D0 U1576 ( .A1(n2256), .A2(port_dest[1]), .ZN(n2253) );
  MUX2D0 U1577 ( .I0(port_dest[0]), .I1(n2257), .S(n2250), .Z(N1449) );
  OAI21D0 U1578 ( .A1(n2249), .A2(n2258), .B(n2251), .ZN(n2257) );
  AOI21D0 U1579 ( .A1(n2259), .A2(n2260), .B(n2255), .ZN(n2258) );
  NR3D0 U1580 ( .A1(n2261), .A2(n2262), .A3(n2263), .ZN(n2255) );
  OAI32D0 U1581 ( .A1(n2264), .A2(n2265), .A3(n2266), .B1(n2267), .B2(n2268), 
        .ZN(n2259) );
  NR2D0 U1582 ( .A1(n2269), .A2(port_dest[0]), .ZN(n2264) );
  INR4D0 U1583 ( .A1(n2263), .B1(n2270), .B2(n2261), .B3(n2262), .ZN(n2249) );
  ND4D0 U1584 ( .A1(n2256), .A2(n2251), .A3(n2252), .A4(n2271), .ZN(N1448) );
  AN4D0 U1585 ( .A1(n2250), .A2(n2260), .A3(n2270), .A4(n2263), .Z(n2271) );
  CKND0 U1586 ( .I(n2254), .ZN(n2260) );
  NR2D0 U1587 ( .A1(n2272), .A2(n2261), .ZN(n2254) );
  IAO21D0 U1588 ( .A1(n2267), .A2(n2268), .B(n2266), .ZN(n2252) );
  AN3D0 U1589 ( .A1(n2273), .A2(n2138), .A3(n2256), .Z(n2266) );
  ND4D0 U1590 ( .A1(n2263), .A2(n2270), .A3(n2274), .A4(n2275), .ZN(n2251) );
  NR3D0 U1591 ( .A1(n2261), .A2(n2262), .A3(n2142), .ZN(n2275) );
  CKND0 U1592 ( .I(n2272), .ZN(n2262) );
  OAI21D0 U1593 ( .A1(port_dest[7]), .A2(n2276), .B(n2277), .ZN(n2272) );
  IND2D0 U1594 ( .A1(n2267), .B1(n2268), .ZN(n2261) );
  OAI21D0 U1595 ( .A1(n2273), .A2(n2138), .B(n2143), .ZN(n2268) );
  IOA21D0 U1596 ( .A1(n2138), .A2(n2273), .B(n2256), .ZN(n2267) );
  IND2D0 U1597 ( .A1(n2278), .B1(n2279), .ZN(n2270) );
  CKND2D0 U1598 ( .A1(n2280), .A2(n2281), .ZN(n2263) );
  NR2D0 U1599 ( .A1(n2265), .A2(n2269), .ZN(n2256) );
  OA21D0 U1600 ( .A1(port_dest[7]), .A2(n2282), .B(n2283), .Z(n2269) );
  AN2D0 U1601 ( .A1(n2282), .A2(port_dest[7]), .Z(n2265) );
  OAI221D0 U1602 ( .A1(port_dest[7]), .A2(n2137), .B1(n2138), .B2(n2284), .C(
        n2285), .ZN(N1366) );
  AOI221D0 U1603 ( .A1(n2278), .A2(n2279), .B1(port_dest[5]), .B2(n2286), .C(
        n2113), .ZN(n2285) );
  AO31D0 U1604 ( .A1(n2287), .A2(n2140), .A3(n2139), .B(port_dest[7]), .Z(
        n2286) );
  CKND2D0 U1605 ( .A1(n2288), .A2(n2280), .ZN(n2139) );
  OAI221D0 U1606 ( .A1(n2289), .A2(n2281), .B1(n2112), .B2(n2290), .C(n2291), 
        .ZN(N1365) );
  AOI31D0 U1607 ( .A1(n2141), .A2(n2140), .A3(n2292), .B(n2113), .ZN(n2291) );
  NR2D0 U1608 ( .A1(n2142), .A2(n2274), .ZN(n2113) );
  IND2D0 U1609 ( .A1(n2279), .B1(n2278), .ZN(n2274) );
  NR2D0 U1610 ( .A1(n2281), .A2(n2280), .ZN(n2278) );
  CKND2D0 U1611 ( .A1(n2293), .A2(n2294), .ZN(n2142) );
  OAI33D0 U1612 ( .A1(n2284), .A2(n2273), .A3(n2138), .B1(n2295), .B2(
        port_dest[7]), .B3(n2282), .ZN(n2292) );
  OAI21D0 U1613 ( .A1(n2283), .A2(port_dest[4]), .B(n2137), .ZN(n2295) );
  CKND2D0 U1614 ( .A1(n2273), .A2(n2287), .ZN(n2137) );
  CKND2D0 U1615 ( .A1(n2287), .A2(n2112), .ZN(n2138) );
  CKND2D0 U1616 ( .A1(n2115), .A2(n2277), .ZN(n2140) );
  CKND2D0 U1617 ( .A1(n2279), .A2(n2288), .ZN(n2141) );
  AOI21D0 U1618 ( .A1(n2296), .A2(n2297), .B(n2298), .ZN(n2279) );
  CKND2D0 U1619 ( .A1(n2288), .A2(n2112), .ZN(n2281) );
  NR2D0 U1620 ( .A1(n2276), .A2(n2277), .ZN(n2288) );
  AOI21D0 U1621 ( .A1(n2296), .A2(n2299), .B(n2300), .ZN(n2277) );
  CKND0 U1622 ( .I(n2115), .ZN(n2276) );
  INR3D0 U1623 ( .A1(n2287), .B1(n2273), .B2(n2143), .ZN(n2115) );
  CKND0 U1624 ( .I(n2284), .ZN(n2143) );
  OAI21D0 U1625 ( .A1(port_dest[11]), .A2(n2301), .B(n2302), .ZN(n2284) );
  NR2D0 U1626 ( .A1(n2303), .A2(n2304), .ZN(n2273) );
  NR2D0 U1627 ( .A1(n2283), .A2(n2282), .ZN(n2287) );
  NR2D0 U1628 ( .A1(n2305), .A2(n2296), .ZN(n2282) );
  AN2D0 U1629 ( .A1(n2306), .A2(n2307), .Z(n2283) );
  CKND0 U1630 ( .I(n2280), .ZN(n2289) );
  AOI31D0 U1631 ( .A1(n2299), .A2(n2296), .A3(n2300), .B(n2308), .ZN(n2280) );
  OAI221D0 U1632 ( .A1(n2309), .A2(n2310), .B1(port_dest[11]), .B2(n2311), .C(
        n2312), .ZN(N1253) );
  NR2D0 U1633 ( .A1(n2299), .A2(port_dest[11]), .ZN(n2309) );
  CKND2D0 U1634 ( .A1(n2313), .A2(n2312), .ZN(N1252) );
  MAOI22D0 U1635 ( .A1(n2296), .A2(n2314), .B1(n2315), .B2(n2294), .ZN(n2312)
         );
  AOI31D0 U1636 ( .A1(n2316), .A2(n2296), .A3(n2311), .B(n2317), .ZN(n2313) );
  OAI31D0 U1637 ( .A1(n2318), .A2(n2307), .A3(n2319), .B(n2320), .ZN(n2316) );
  OAI21D0 U1638 ( .A1(n2315), .A2(n2294), .B(n2321), .ZN(N1251) );
  MUX2ND0 U1639 ( .I0(n2322), .I1(port_dest[8]), .S(port_dest[11]), .ZN(n2321)
         );
  NR2D0 U1640 ( .A1(n2314), .A2(n2323), .ZN(n2322) );
  AOI21D0 U1641 ( .A1(n2324), .A2(n2325), .B(n2326), .ZN(n2323) );
  OAI32D0 U1642 ( .A1(n2327), .A2(n2319), .A3(n2328), .B1(n2301), .B2(n2329), 
        .ZN(n2324) );
  NR2D0 U1643 ( .A1(n2307), .A2(port_dest[8]), .ZN(n2327) );
  ND3D0 U1644 ( .A1(n2298), .A2(n2296), .A3(n2297), .ZN(n2294) );
  CKND0 U1645 ( .I(n2330), .ZN(n2297) );
  CKND0 U1646 ( .I(n2293), .ZN(n2315) );
  ND4D0 U1647 ( .A1(n2311), .A2(n2304), .A3(n2331), .A4(n2320), .ZN(N1250) );
  IAO21D0 U1648 ( .A1(n2301), .A2(n2329), .B(n2328), .ZN(n2320) );
  NR3D0 U1649 ( .A1(n2319), .A2(n2307), .A3(n2303), .ZN(n2328) );
  CKND0 U1650 ( .I(n2305), .ZN(n2319) );
  NR2D0 U1651 ( .A1(n2293), .A2(n2314), .ZN(n2331) );
  NR2D0 U1652 ( .A1(n2298), .A2(n2330), .ZN(n2314) );
  ND3D0 U1653 ( .A1(n2300), .A2(n2308), .A3(n2299), .ZN(n2330) );
  CKND0 U1654 ( .I(n2332), .ZN(n2300) );
  OAI21D0 U1655 ( .A1(n2333), .A2(n2334), .B(n2335), .ZN(n2298) );
  NR2D0 U1656 ( .A1(n2336), .A2(n2337), .ZN(n2293) );
  NR2D0 U1657 ( .A1(n2306), .A2(n2307), .ZN(n2304) );
  CKND0 U1658 ( .I(n2338), .ZN(n2307) );
  CKND2D0 U1659 ( .A1(n2296), .A2(n2305), .ZN(n2306) );
  INR2D0 U1660 ( .A1(n2325), .B1(n2326), .ZN(n2311) );
  INR3D0 U1661 ( .A1(n2299), .B1(n2332), .B2(n2308), .ZN(n2326) );
  CKND2D0 U1662 ( .A1(n2333), .A2(n2334), .ZN(n2308) );
  CKND2D0 U1663 ( .A1(n2332), .A2(n2299), .ZN(n2325) );
  NR2D0 U1664 ( .A1(n2301), .A2(n2302), .ZN(n2299) );
  CKND0 U1665 ( .I(n2329), .ZN(n2302) );
  OAI21D0 U1666 ( .A1(port_dest[15]), .A2(n2339), .B(n2340), .ZN(n2329) );
  ND3D0 U1667 ( .A1(n2305), .A2(n2338), .A3(n2303), .ZN(n2301) );
  OAI21D0 U1668 ( .A1(n2341), .A2(n2342), .B(n2343), .ZN(n2303) );
  CKND2D0 U1669 ( .A1(n2341), .A2(n2342), .ZN(n2338) );
  CKND2D0 U1670 ( .A1(n2344), .A2(port_dest[15]), .ZN(n2305) );
  AOI21D0 U1671 ( .A1(n2345), .A2(n2346), .B(n2347), .ZN(n2332) );
  OAI211D0 U1672 ( .A1(port_dest[15]), .A2(n2348), .B(n2349), .C(n2350), .ZN(
        N1139) );
  NR4D0 U1673 ( .A1(n2351), .A2(n2352), .A3(n2353), .A4(n2354), .ZN(n2348) );
  AN2D0 U1674 ( .A1(port_dest[14]), .A2(n2346), .Z(n2354) );
  OAI221D0 U1675 ( .A1(n2355), .A2(n2356), .B1(port_dest[15]), .B2(n2357), .C(
        n2349), .ZN(N1138) );
  AOI31D0 U1676 ( .A1(n2358), .A2(n2359), .A3(n2360), .B(port_dest[15]), .ZN(
        n2355) );
  CKND2D0 U1677 ( .A1(n2361), .A2(n2349), .ZN(N1137) );
  IND2D0 U1678 ( .A1(n2336), .B1(n2337), .ZN(n2349) );
  NR3D0 U1679 ( .A1(n2335), .A2(n2333), .A3(n2334), .ZN(n2337) );
  CKND2D0 U1680 ( .A1(n2362), .A2(n2345), .ZN(n2334) );
  MUX2ND0 U1681 ( .I0(n2363), .I1(port_dest[12]), .S(port_dest[15]), .ZN(n2361) );
  NR2D0 U1682 ( .A1(n2351), .A2(n2364), .ZN(n2363) );
  AOI21D0 U1683 ( .A1(n2365), .A2(n2359), .B(n2353), .ZN(n2364) );
  OAI22D0 U1684 ( .A1(n2339), .A2(n2366), .B1(n2344), .B2(n2367), .ZN(n2365)
         );
  AOI21D0 U1685 ( .A1(port_dest[12]), .A2(n2368), .B(n2341), .ZN(n2367) );
  IND4D0 U1686 ( .A1(n2341), .B1(n2369), .B2(n2336), .B3(n2359), .ZN(N1136) );
  CKND0 U1687 ( .I(n2352), .ZN(n2359) );
  NR2D0 U1688 ( .A1(n2347), .A2(n2370), .ZN(n2352) );
  OAI31D0 U1689 ( .A1(n2182), .A2(n2371), .A3(n2372), .B(n2373), .ZN(n2336) );
  INR3D0 U1690 ( .A1(n2357), .B1(n2353), .B2(n2342), .ZN(n2369) );
  OR2D0 U1691 ( .A1(n2344), .A2(port_dest[15]), .Z(n2342) );
  CKND0 U1692 ( .I(n2358), .ZN(n2353) );
  CKND2D0 U1693 ( .A1(n2333), .A2(n2362), .ZN(n2358) );
  CKND0 U1694 ( .I(n2374), .ZN(n2333) );
  AOI221D0 U1695 ( .A1(n2360), .A2(n2343), .B1(n2375), .B2(n2340), .C(n2351), 
        .ZN(n2357) );
  AN3D0 U1696 ( .A1(n2362), .A2(n2374), .A3(n2335), .Z(n2351) );
  OA31D0 U1697 ( .A1(n2182), .A2(n2371), .A3(n2376), .B(n2377), .Z(n2335) );
  OAI21D0 U1698 ( .A1(n2376), .A2(n2182), .B(n2371), .ZN(n2374) );
  AN2D0 U1699 ( .A1(n2347), .A2(n2346), .Z(n2362) );
  CKND0 U1700 ( .I(n2370), .ZN(n2346) );
  CKND2D0 U1701 ( .A1(n2375), .A2(n2366), .ZN(n2370) );
  CKND2D0 U1702 ( .A1(n2376), .A2(n2182), .ZN(n2347) );
  CKND0 U1703 ( .I(n2366), .ZN(n2340) );
  OAI21D0 U1704 ( .A1(port_dest[19]), .A2(n2378), .B(n2379), .ZN(n2366) );
  CKND0 U1705 ( .I(n2339), .ZN(n2375) );
  CKND2D0 U1706 ( .A1(n2360), .A2(n2368), .ZN(n2339) );
  CKND0 U1707 ( .I(n2368), .ZN(n2343) );
  OAI21D0 U1708 ( .A1(port_dest[19]), .A2(n2380), .B(n2381), .ZN(n2368) );
  NR2D0 U1709 ( .A1(n2341), .A2(n2344), .ZN(n2360) );
  NR2D0 U1710 ( .A1(n2382), .A2(n2383), .ZN(n2344) );
  AOI21D0 U1711 ( .A1(n2383), .A2(n2382), .B(n2384), .ZN(n2341) );
  OAI221D0 U1712 ( .A1(port_dest[19]), .A2(n2183), .B1(n2385), .B2(n2182), .C(
        n2386), .ZN(N1025) );
  CKND0 U1713 ( .I(port_dest[18]), .ZN(n2385) );
  OAI31D0 U1714 ( .A1(n2372), .A2(n2371), .A3(n2373), .B(n2387), .ZN(n2183) );
  OAI31D0 U1715 ( .A1(n2182), .A2(n2376), .A3(n2388), .B(n2389), .ZN(N1024) );
  MUX2ND0 U1716 ( .I0(n2390), .I1(port_dest[16]), .S(port_dest[19]), .ZN(n2389) );
  AOI21D0 U1717 ( .A1(n2387), .A2(n2372), .B(n2391), .ZN(n2390) );
  AOI22D0 U1718 ( .A1(n2392), .A2(n2382), .B1(n2379), .B2(n2393), .ZN(n2391)
         );
  OAI21D0 U1719 ( .A1(n2381), .A2(n2394), .B(n2384), .ZN(n2392) );
  OR2D0 U1720 ( .A1(n2376), .A2(n2377), .Z(n2372) );
  AOI21D0 U1721 ( .A1(n2373), .A2(n2395), .B(n2371), .ZN(n2388) );
  NR2D0 U1722 ( .A1(n2396), .A2(n2397), .ZN(n2371) );
  CKND0 U1723 ( .I(n2377), .ZN(n2395) );
  AOI21D0 U1724 ( .A1(n2396), .A2(n2397), .B(n2204), .ZN(n2377) );
  AN2D0 U1725 ( .A1(n2185), .A2(n2193), .Z(n2373) );
  ND3D0 U1726 ( .A1(n2204), .A2(n2396), .A3(n2397), .ZN(n2193) );
  NR2D0 U1727 ( .A1(n2198), .A2(port_dest[23]), .ZN(n2397) );
  CKND2D0 U1728 ( .A1(n2154), .A2(n2203), .ZN(n2198) );
  CKND0 U1729 ( .I(n2191), .ZN(n2396) );
  NR2D0 U1730 ( .A1(n2219), .A2(n2398), .ZN(n2191) );
  CKND2D0 U1731 ( .A1(n2223), .A2(n2218), .ZN(n2204) );
  IAO21D0 U1732 ( .A1(n2223), .A2(n2218), .B(n2213), .ZN(n2185) );
  IND2D0 U1733 ( .A1(n2226), .B1(n2229), .ZN(n2213) );
  ND3D0 U1734 ( .A1(n2244), .A2(n2232), .A3(n2399), .ZN(n2229) );
  ND4D0 U1735 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2226) );
  AOI33D0 U1736 ( .A1(port_dest[0]), .A2(n2404), .A3(port_dest[2]), .B1(
        port_dest[8]), .B2(n2317), .B3(port_dest[10]), .ZN(n2403) );
  AOI33D0 U1737 ( .A1(port_dest[20]), .A2(port_dest[21]), .A3(n2405), .B1(
        port_dest[24]), .B2(port_dest[25]), .B3(n2210), .ZN(n2402) );
  AOI33D0 U1738 ( .A1(port_dest[28]), .A2(port_dest[29]), .A3(n2173), .B1(
        port_dest[4]), .B2(port_dest[5]), .B3(n2114), .ZN(n2401) );
  AOI33D0 U1739 ( .A1(port_dest[12]), .A2(port_dest[13]), .A3(n2406), .B1(
        port_dest[16]), .B2(port_dest[17]), .B3(n2407), .ZN(n2400) );
  CKND2D0 U1740 ( .A1(n2398), .A2(n2219), .ZN(n2218) );
  CKND0 U1741 ( .I(n2225), .ZN(n2219) );
  NR2D0 U1742 ( .A1(n2244), .A2(n2399), .ZN(n2225) );
  NR2D0 U1743 ( .A1(n2206), .A2(n2224), .ZN(n2398) );
  AOI21D0 U1744 ( .A1(n2244), .A2(n2399), .B(n2232), .ZN(n2223) );
  ND4D0 U1745 ( .A1(n2408), .A2(n2409), .A3(n2410), .A4(n2411), .ZN(n2232) );
  AOI33D0 U1746 ( .A1(n2317), .A2(n2412), .A3(port_dest[10]), .B1(n2404), .B2(
        n2413), .B3(port_dest[2]), .ZN(n2411) );
  AOI33D0 U1747 ( .A1(port_dest[17]), .A2(n2394), .A3(n2407), .B1(
        port_dest[13]), .B2(n2414), .B3(n2406), .ZN(n2410) );
  AOI33D0 U1748 ( .A1(port_dest[5]), .A2(n2290), .A3(n2114), .B1(port_dest[29]), .B2(n2415), .B3(n2173), .ZN(n2409) );
  AOI33D0 U1749 ( .A1(port_dest[25]), .A2(n2416), .A3(n2210), .B1(
        port_dest[21]), .B2(n2417), .B3(n2405), .ZN(n2408) );
  NR2D0 U1750 ( .A1(n2171), .A2(n2239), .ZN(n2399) );
  ND4D0 U1751 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(n2244) );
  AOI33D0 U1752 ( .A1(port_dest[8]), .A2(n2422), .A3(port_dest[10]), .B1(
        port_dest[0]), .B2(n2423), .B3(port_dest[2]), .ZN(n2421) );
  AOI33D0 U1753 ( .A1(port_dest[20]), .A2(n2176), .A3(n2405), .B1(
        port_dest[24]), .B2(n2215), .B3(n2210), .ZN(n2420) );
  AOI33D0 U1754 ( .A1(port_dest[28]), .A2(n2168), .A3(n2173), .B1(port_dest[4]), .B2(n2424), .B3(n2114), .ZN(n2419) );
  AOI33D0 U1755 ( .A1(port_dest[12]), .A2(n2356), .A3(n2406), .B1(
        port_dest[16]), .B2(n2425), .B3(n2407), .ZN(n2418) );
  AOI21D0 U1756 ( .A1(n2426), .A2(n2154), .B(n2203), .ZN(n2376) );
  CKND2D0 U1757 ( .A1(n2224), .A2(n2206), .ZN(n2203) );
  CKND0 U1758 ( .I(n2211), .ZN(n2206) );
  INR2D0 U1759 ( .A1(n2216), .B1(n2217), .ZN(n2211) );
  NR2D0 U1760 ( .A1(n2427), .A2(n2428), .ZN(n2216) );
  CKND0 U1761 ( .I(n2220), .ZN(n2224) );
  CKND2D0 U1762 ( .A1(n2239), .A2(n2171), .ZN(n2220) );
  CKND2D0 U1763 ( .A1(n2165), .A2(n2237), .ZN(n2171) );
  CKND0 U1764 ( .I(n2235), .ZN(n2239) );
  ND4D0 U1765 ( .A1(n2429), .A2(n2430), .A3(n2431), .A4(n2432), .ZN(n2235) );
  AOI33D0 U1766 ( .A1(n2422), .A2(n2412), .A3(port_dest[10]), .B1(n2423), .B2(
        n2413), .B3(port_dest[2]), .ZN(n2432) );
  AOI33D0 U1767 ( .A1(n2417), .A2(n2176), .A3(n2405), .B1(n2416), .B2(n2215), 
        .B3(n2210), .ZN(n2431) );
  NR2D0 U1768 ( .A1(n2205), .A2(n2433), .ZN(n2210) );
  CKND0 U1769 ( .I(port_dest[26]), .ZN(n2205) );
  CKND0 U1770 ( .I(n2152), .ZN(n2405) );
  CKND2D0 U1771 ( .A1(port_dest[22]), .A2(port_dest[23]), .ZN(n2152) );
  AOI33D0 U1772 ( .A1(n2415), .A2(n2168), .A3(n2173), .B1(n2290), .B2(n2424), 
        .B3(n2114), .ZN(n2430) );
  AN2D0 U1773 ( .A1(port_dest[6]), .A2(port_dest[7]), .Z(n2114) );
  NR2D0 U1774 ( .A1(n2170), .A2(n2434), .ZN(n2173) );
  CKND0 U1775 ( .I(port_dest[30]), .ZN(n2170) );
  AOI33D0 U1776 ( .A1(n2414), .A2(n2356), .A3(n2406), .B1(n2394), .B2(n2425), 
        .B3(n2407), .ZN(n2429) );
  CKND0 U1777 ( .I(n2386), .ZN(n2407) );
  CKND2D0 U1778 ( .A1(port_dest[18]), .A2(port_dest[19]), .ZN(n2386) );
  CKND0 U1779 ( .I(n2350), .ZN(n2406) );
  CKND2D0 U1780 ( .A1(port_dest[14]), .A2(port_dest[15]), .ZN(n2350) );
  INR2D0 U1781 ( .A1(n2187), .B1(n2186), .ZN(n2154) );
  CKND2D0 U1782 ( .A1(n2387), .A2(n2383), .ZN(n2182) );
  NR2D0 U1783 ( .A1(n2378), .A2(n2379), .ZN(n2387) );
  IAO21D0 U1784 ( .A1(port_dest[23]), .A2(n2186), .B(n2187), .ZN(n2379) );
  OAI21D0 U1785 ( .A1(n2428), .A2(n2217), .B(n2427), .ZN(n2187) );
  NR2D0 U1786 ( .A1(n2237), .A2(n2165), .ZN(n2427) );
  NR2D0 U1787 ( .A1(n2240), .A2(port_dest[31]), .ZN(n2165) );
  CKND2D0 U1788 ( .A1(n2163), .A2(n2167), .ZN(n2240) );
  ND4D0 U1789 ( .A1(n2435), .A2(n2436), .A3(n2437), .A4(n2438), .ZN(n2237) );
  AOI33D0 U1790 ( .A1(port_dest[17]), .A2(n2439), .A3(port_dest[16]), .B1(
        port_dest[13]), .B2(n2440), .B3(port_dest[12]), .ZN(n2438) );
  AOI33D0 U1791 ( .A1(port_dest[5]), .A2(n2441), .A3(port_dest[4]), .B1(
        port_dest[25]), .B2(n2442), .B3(port_dest[24]), .ZN(n2437) );
  AOI33D0 U1792 ( .A1(port_dest[29]), .A2(n2443), .A3(port_dest[28]), .B1(
        port_dest[21]), .B2(n2444), .B3(port_dest[20]), .ZN(n2436) );
  AOI33D0 U1793 ( .A1(n2404), .A2(n2445), .A3(port_dest[0]), .B1(n2317), .B2(
        n2310), .B3(port_dest[8]), .ZN(n2435) );
  CKND2D0 U1794 ( .A1(n2181), .A2(n2201), .ZN(n2186) );
  CKND0 U1795 ( .I(n2393), .ZN(n2378) );
  NR2D0 U1796 ( .A1(n2380), .A2(n2381), .ZN(n2393) );
  AOI21D0 U1797 ( .A1(n2426), .A2(n2181), .B(n2201), .ZN(n2381) );
  CKND2D0 U1798 ( .A1(n2428), .A2(n2217), .ZN(n2201) );
  CKND2D0 U1799 ( .A1(n2221), .A2(n2433), .ZN(n2217) );
  AOI21D0 U1800 ( .A1(port_dest[31]), .A2(n2241), .B(n2446), .ZN(n2221) );
  AOI21D0 U1801 ( .A1(n2434), .A2(n2163), .B(n2167), .ZN(n2428) );
  ND4D0 U1802 ( .A1(n2447), .A2(n2448), .A3(n2449), .A4(n2450), .ZN(n2167) );
  AOI33D0 U1803 ( .A1(n2439), .A2(n2394), .A3(port_dest[17]), .B1(n2440), .B2(
        n2414), .B3(port_dest[13]), .ZN(n2450) );
  AOI33D0 U1804 ( .A1(n2441), .A2(n2290), .A3(port_dest[5]), .B1(n2442), .B2(
        n2416), .B3(port_dest[25]), .ZN(n2449) );
  AOI33D0 U1805 ( .A1(n2443), .A2(n2415), .A3(port_dest[29]), .B1(n2444), .B2(
        n2417), .B3(port_dest[21]), .ZN(n2448) );
  AOI33D0 U1806 ( .A1(n2413), .A2(n2445), .A3(n2404), .B1(n2310), .B2(n2412), 
        .B3(n2317), .ZN(n2447) );
  NR2D0 U1807 ( .A1(n2318), .A2(n2296), .ZN(n2317) );
  CKND0 U1808 ( .I(port_dest[9]), .ZN(n2318) );
  CKND0 U1809 ( .I(n2245), .ZN(n2404) );
  CKND2D0 U1810 ( .A1(port_dest[3]), .A2(port_dest[1]), .ZN(n2245) );
  NR2D0 U1811 ( .A1(n2241), .A2(n2243), .ZN(n2163) );
  CKND0 U1812 ( .I(n2451), .ZN(n2243) );
  CKND0 U1813 ( .I(n2452), .ZN(n2241) );
  NR2D0 U1814 ( .A1(n2202), .A2(n2200), .ZN(n2181) );
  CKND2D0 U1815 ( .A1(n2384), .A2(n2382), .ZN(n2380) );
  CKND2D0 U1816 ( .A1(n2200), .A2(port_dest[23]), .ZN(n2382) );
  OAI21D0 U1817 ( .A1(port_dest[23]), .A2(n2200), .B(n2202), .ZN(n2384) );
  AN2D0 U1818 ( .A1(n2446), .A2(n2453), .Z(n2202) );
  OAI21D0 U1819 ( .A1(n2434), .A2(n2452), .B(n2433), .ZN(n2453) );
  AOI21D0 U1820 ( .A1(n2434), .A2(n2452), .B(n2451), .ZN(n2446) );
  ND4D0 U1821 ( .A1(n2454), .A2(n2455), .A3(n2456), .A4(n2457), .ZN(n2451) );
  AOI33D0 U1822 ( .A1(n2439), .A2(n2425), .A3(port_dest[16]), .B1(n2440), .B2(
        n2356), .B3(port_dest[12]), .ZN(n2457) );
  AOI33D0 U1823 ( .A1(n2422), .A2(n2310), .A3(port_dest[8]), .B1(n2441), .B2(
        n2424), .B3(port_dest[4]), .ZN(n2456) );
  AOI33D0 U1824 ( .A1(n2423), .A2(n2445), .A3(port_dest[0]), .B1(n2442), .B2(
        n2215), .B3(port_dest[24]), .ZN(n2455) );
  AOI33D0 U1825 ( .A1(n2443), .A2(n2168), .A3(port_dest[28]), .B1(n2444), .B2(
        n2176), .B3(port_dest[20]), .ZN(n2454) );
  NR3D0 U1826 ( .A1(n2434), .A2(n2433), .A3(n2452), .ZN(n2200) );
  ND4D0 U1827 ( .A1(n2458), .A2(n2459), .A3(n2460), .A4(n2461), .ZN(n2452) );
  AOI33D0 U1828 ( .A1(n2394), .A2(n2425), .A3(n2439), .B1(n2414), .B2(n2356), 
        .B3(n2440), .ZN(n2461) );
  NR2D0 U1829 ( .A1(n2345), .A2(port_dest[14]), .ZN(n2440) );
  CKND0 U1830 ( .I(port_dest[15]), .ZN(n2345) );
  CKND0 U1831 ( .I(port_dest[13]), .ZN(n2356) );
  CKND0 U1832 ( .I(port_dest[12]), .ZN(n2414) );
  NR2D0 U1833 ( .A1(n2383), .A2(port_dest[18]), .ZN(n2439) );
  CKND0 U1834 ( .I(port_dest[19]), .ZN(n2383) );
  CKND0 U1835 ( .I(port_dest[17]), .ZN(n2425) );
  CKND0 U1836 ( .I(port_dest[16]), .ZN(n2394) );
  AOI33D0 U1837 ( .A1(n2310), .A2(n2412), .A3(n2422), .B1(n2290), .B2(n2424), 
        .B3(n2441), .ZN(n2460) );
  NR2D0 U1838 ( .A1(n2112), .A2(port_dest[6]), .ZN(n2441) );
  CKND0 U1839 ( .I(port_dest[7]), .ZN(n2112) );
  CKND0 U1840 ( .I(port_dest[5]), .ZN(n2424) );
  CKND0 U1841 ( .I(port_dest[4]), .ZN(n2290) );
  NR2D0 U1842 ( .A1(n2296), .A2(port_dest[9]), .ZN(n2422) );
  CKND0 U1843 ( .I(port_dest[11]), .ZN(n2296) );
  CKND0 U1844 ( .I(port_dest[8]), .ZN(n2412) );
  CKND0 U1845 ( .I(port_dest[10]), .ZN(n2310) );
  AOI33D0 U1846 ( .A1(n2413), .A2(n2445), .A3(n2423), .B1(n2416), .B2(n2215), 
        .B3(n2442), .ZN(n2459) );
  NR2D0 U1847 ( .A1(n2433), .A2(port_dest[26]), .ZN(n2442) );
  CKND0 U1848 ( .I(port_dest[25]), .ZN(n2215) );
  CKND0 U1849 ( .I(port_dest[24]), .ZN(n2416) );
  NR2D0 U1850 ( .A1(n2250), .A2(port_dest[1]), .ZN(n2423) );
  CKND0 U1851 ( .I(port_dest[3]), .ZN(n2250) );
  CKND0 U1852 ( .I(port_dest[2]), .ZN(n2445) );
  CKND0 U1853 ( .I(port_dest[0]), .ZN(n2413) );
  AOI33D0 U1854 ( .A1(n2415), .A2(n2168), .A3(n2443), .B1(n2417), .B2(n2176), 
        .B3(n2444), .ZN(n2458) );
  NR2D0 U1855 ( .A1(n2426), .A2(port_dest[22]), .ZN(n2444) );
  CKND0 U1856 ( .I(port_dest[23]), .ZN(n2426) );
  CKND0 U1857 ( .I(port_dest[21]), .ZN(n2176) );
  CKND0 U1858 ( .I(port_dest[20]), .ZN(n2417) );
  NR2D0 U1859 ( .A1(n2434), .A2(port_dest[30]), .ZN(n2443) );
  CKND0 U1860 ( .I(port_dest[29]), .ZN(n2168) );
  CKND0 U1861 ( .I(port_dest[28]), .ZN(n2415) );
  CKND0 U1862 ( .I(port_dest[27]), .ZN(n2433) );
  CKND0 U1863 ( .I(port_dest[31]), .ZN(n2434) );
endmodule

