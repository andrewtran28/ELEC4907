
module routing_engine_CLOCKED ( port_dest, clk, rst, control, done );
  input [31:0] port_dest;
  output [19:0] control;
  input clk, rst;
  output done;
  wire   \dst[0][2] , \dst[0][1] , \dst[0][0] , \dst[1][2] , \dst[1][1] ,
         \dst[1][0] , \dst[2][2] , \dst[2][1] , \dst[2][0] , \dst[3][2] ,
         \dst[3][0] , \dst[4][2] , \dst[4][1] , \dst[4][0] , \dst[5][2] ,
         \dst[5][1] , \dst[5][0] , \dst[6][2] , \dst[6][1] , \dst[6][0] ,
         \dst[7][1] , \dst[7][0] , \stage_1_output[0][1] ,
         \stage_1_output[0][2] , \stage_1_output[1][2] ,
         \stage_1_output[2][1] , \stage_1_output[2][2] ,
         \stage_1_output[3][2] , \stage_1_output[4][1] , N1614, N1615, N1616,
         N1618, n1, n2, n11, n13, n277, n386, n388, n397, n398, n400, n401,
         n403, n41, n370, n371, n375, n376, n6, n7, n8, n14, n17, n18, n19,
         n20, n46, \control[19] , n357, n358, n359, n360, n361, n362, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041;
  assign control[13] = \control[19] ;
  assign control[15] = \control[19] ;
  assign control[19] = \control[19] ;

  DFD1 \stage_1_output_reg[6][1]  ( .D(N1618), .CP(clk), .QN(n1041) );
  EDFQD1 \dst_reg[2][0]  ( .D(n2), .E(n41), .CP(clk), .Q(\dst[2][0] ) );
  EDFQD1 \dst_reg[4][0]  ( .D(n1), .E(n375), .CP(clk), .Q(\dst[4][0] ) );
  EDFQD1 \dst_reg[4][2]  ( .D(n46), .E(n375), .CP(clk), .Q(\dst[4][2] ) );
  EDFQD1 \dst_reg[2][2]  ( .D(n362), .E(n41), .CP(clk), .Q(\dst[2][2] ) );
  EDFQD1 \dst_reg[2][1]  ( .D(n376), .E(n41), .CP(clk), .Q(\dst[2][1] ) );
  DFKCNQD1 \stage_1_output_reg[4][1]  ( .CN(done), .D(n401), .CP(clk), .Q(
        \stage_1_output[4][1] ) );
  DFQD1 \dst_reg[0][0]  ( .D(n403), .CP(clk), .Q(\dst[0][0] ) );
  DFQD1 \dst_reg[1][1]  ( .D(n401), .CP(clk), .Q(\dst[1][1] ) );
  DFQD1 \dst_reg[1][0]  ( .D(n400), .CP(clk), .Q(\dst[1][0] ) );
  DFQD1 \dst_reg[3][2]  ( .D(n13), .CP(clk), .Q(\dst[3][2] ) );
  DFQD1 \dst_reg[1][2]  ( .D(n371), .CP(clk), .Q(\dst[1][2] ) );
  DFQD1 \dst_reg[6][2]  ( .D(n19), .CP(clk), .Q(\dst[6][2] ) );
  DFQD1 \dst_reg[7][0]  ( .D(n386), .CP(clk), .Q(\dst[7][0] ) );
  DFQD1 \dst_reg[0][1]  ( .D(n17), .CP(clk), .Q(\dst[0][1] ) );
  DFQD1 \dst_reg[0][2]  ( .D(n20), .CP(clk), .Q(\dst[0][2] ) );
  DFQD1 \dst_reg[3][0]  ( .D(n397), .CP(clk), .Q(\dst[3][0] ) );
  DFQD1 \dst_reg[6][0]  ( .D(n388), .CP(clk), .Q(\dst[6][0] ) );
  DFQD1 \dst_reg[5][1]  ( .D(n358), .CP(clk), .Q(\dst[5][1] ) );
  DFQD1 \dst_reg[5][0]  ( .D(n359), .CP(clk), .Q(\dst[5][0] ) );
  DFQD1 \dst_reg[5][2]  ( .D(n360), .CP(clk), .Q(\dst[5][2] ) );
  DFQD1 \dst_reg[7][1]  ( .D(n361), .CP(clk), .Q(\dst[7][1] ) );
  DFXQD1 \stage_1_output_reg[0][2]  ( .DB(n400), .DA(n403), .SA(done), .CP(clk), .Q(\stage_1_output[0][2] ) );
  DFXQD1 \stage_1_output_reg[1][2]  ( .DB(n397), .DA(n398), .SA(n370), .CP(clk), .Q(\stage_1_output[1][2] ) );
  DFQD1 \stage_1_output_reg[0][1]  ( .D(n17), .CP(clk), .Q(
        \stage_1_output[0][1] ) );
  DFQD1 \stage_1_output_reg[2][1]  ( .D(N1615), .CP(clk), .Q(
        \stage_1_output[2][1] ) );
  DFQD1 \dst_reg[6][1]  ( .D(n18), .CP(clk), .Q(\dst[6][1] ) );
  DFQD1 \stage_1_output_reg[2][2]  ( .D(N1614), .CP(clk), .Q(
        \stage_1_output[2][2] ) );
  DFQD1 \stage_1_output_reg[3][2]  ( .D(N1616), .CP(clk), .Q(
        \stage_1_output[3][2] ) );
  EDFQD1 \dst_reg[4][1]  ( .D(n277), .E(n375), .CP(clk), .Q(\dst[4][1] ) );
  DFQD1 \stage_0_sw_ctl_reg[1]  ( .D(n14), .CP(clk), .Q(control[18]) );
  DFQD1 \stage_0_sw_ctl_reg[2]  ( .D(n7), .CP(clk), .Q(control[17]) );
  DFQD1 \stage_1_sw_ctl_reg[3]  ( .D(n357), .CP(clk), .Q(control[12]) );
  DFQD1 \stage_1_sw_ctl_reg[1]  ( .D(n6), .CP(clk), .Q(control[14]) );
  DFQD1 \stage_0_sw_ctl_reg[3]  ( .D(n8), .CP(clk), .Q(control[16]) );
  DFKCNQD1 \stage_1_output_reg[4][0]  ( .CN(done), .D(n371), .CP(clk), .Q(
        control[9]) );
  DFQD1 \stage_1_output_reg[0][0]  ( .D(n20), .CP(clk), .Q(control[11]) );
  DFXQD1 \stage_1_output_reg[5][0]  ( .DB(n11), .DA(n13), .SA(n370), .CP(clk), 
        .Q(control[8]) );
  DFXQD1 \stage_1_output_reg[1][0]  ( .DB(n13), .DA(n11), .SA(n370), .CP(clk), 
        .Q(control[10]) );
  MUX2ND1 U3 ( .I0(n772), .I1(n771), .S(control[6]), .ZN(control[0]) );
  MUX2ND1 U4 ( .I0(n770), .I1(n769), .S(control[7]), .ZN(control[2]) );
  MUX2ND1 U5 ( .I0(n769), .I1(n770), .S(control[7]), .ZN(control[3]) );
  CKMUX2D1 U6 ( .I0(\stage_1_output[0][1] ), .I1(\stage_1_output[2][1] ), .S(
        control[11]), .Z(control[7]) );
  MUX2ND1 U7 ( .I0(n771), .I1(n772), .S(control[6]), .ZN(control[1]) );
  MUX2ND1 U8 ( .I0(n1041), .I1(n768), .S(control[9]), .ZN(control[4]) );
  CKMUX2D1 U9 ( .I0(\stage_1_output[2][1] ), .I1(\stage_1_output[0][1] ), .S(
        control[11]), .Z(control[6]) );
  MUX2ND1 U10 ( .I0(n768), .I1(n1041), .S(control[9]), .ZN(control[5]) );
  TIEH U11 ( .Z(done) );
  TIEL U12 ( .ZN(\control[19] ) );
  MUX2D0 U13 ( .I0(\dst[0][0] ), .I1(n713), .S(n714), .Z(n403) );
  OAI32D0 U14 ( .A1(n715), .A2(n716), .A3(n717), .B1(n718), .B2(n719), .ZN(
        n713) );
  OAI21D0 U15 ( .A1(n720), .A2(n721), .B(n722), .ZN(n715) );
  MUX2D0 U16 ( .I0(\dst[1][1] ), .I1(n723), .S(n724), .Z(n401) );
  OAI211D0 U17 ( .A1(n725), .A2(n726), .B(n727), .C(n728), .ZN(n723) );
  MUX2ND0 U18 ( .I0(port_dest[25]), .I1(n729), .S(n730), .ZN(n728) );
  CKND0 U19 ( .I(n731), .ZN(n725) );
  MUX2D0 U20 ( .I0(\dst[1][0] ), .I1(n732), .S(n724), .Z(n400) );
  OAI32D0 U21 ( .A1(n733), .A2(n729), .A3(n734), .B1(n730), .B2(n735), .ZN(
        n732) );
  MUX2D0 U22 ( .I0(\dst[2][0] ), .I1(n2), .S(n41), .Z(n398) );
  MUX3D0 U23 ( .I0(port_dest[16]), .I1(n736), .I2(\dst[3][0] ), .S0(n737), 
        .S1(n738), .Z(n397) );
  OA211D0 U24 ( .A1(n739), .A2(n740), .B(n741), .C(n742), .Z(n736) );
  CKND0 U25 ( .I(n743), .ZN(n740) );
  MUX2D0 U26 ( .I0(n744), .I1(port_dest[20]), .S(port_dest[23]), .Z(n2) );
  AOI211D0 U27 ( .A1(n745), .A2(n746), .B(n747), .C(n748), .ZN(n744) );
  CKND2D0 U28 ( .A1(n749), .A2(n733), .ZN(n746) );
  CKND0 U29 ( .I(n370), .ZN(n14) );
  OAI221D0 U30 ( .A1(n750), .A2(n751), .B1(n752), .B2(n753), .C(n754), .ZN(
        n370) );
  AN2D0 U31 ( .A1(n755), .A2(n756), .Z(n754) );
  OAI221D0 U32 ( .A1(port_dest[19]), .A2(n741), .B1(n757), .B2(n758), .C(n759), 
        .ZN(n13) );
  AOI221D0 U33 ( .A1(\dst[3][2] ), .A2(n738), .B1(n760), .B2(n761), .C(n762), 
        .ZN(n759) );
  AN4D0 U34 ( .A1(n763), .A2(n761), .A3(n741), .A4(n758), .Z(n738) );
  CKND0 U35 ( .I(n760), .ZN(n763) );
  CKND2D0 U36 ( .A1(n764), .A2(n765), .ZN(n741) );
  OAI21D0 U37 ( .A1(n760), .A2(n766), .B(n767), .ZN(n765) );
  CKND0 U38 ( .I(\stage_1_output[4][1] ), .ZN(n768) );
  MUX2ND0 U39 ( .I0(\stage_1_output[0][2] ), .I1(\stage_1_output[2][2] ), .S(
        control[11]), .ZN(n769) );
  MUX2ND0 U40 ( .I0(\stage_1_output[1][2] ), .I1(\stage_1_output[3][2] ), .S(
        control[10]), .ZN(n770) );
  MUX2ND0 U41 ( .I0(\stage_1_output[2][2] ), .I1(\stage_1_output[0][2] ), .S(
        control[11]), .ZN(n771) );
  MUX2ND0 U42 ( .I0(\stage_1_output[3][2] ), .I1(\stage_1_output[1][2] ), .S(
        control[10]), .ZN(n772) );
  MUX3ND0 U43 ( .I0(n773), .I1(n774), .I2(n775), .S0(n7), .S1(n357), .ZN(N1618) );
  CKXOR2D0 U44 ( .A1(n776), .A2(n371), .Z(n357) );
  OA32D0 U45 ( .A1(n777), .A2(n778), .A3(n779), .B1(\dst[1][2] ), .B2(n724), 
        .Z(n371) );
  ND3D0 U46 ( .A1(n780), .A2(n731), .A3(n781), .ZN(n724) );
  AOI211D0 U47 ( .A1(n782), .A2(n783), .B(n784), .C(n729), .ZN(n781) );
  NR3D0 U48 ( .A1(n749), .A2(n785), .A3(n786), .ZN(n729) );
  CKND2D0 U49 ( .A1(n787), .A2(n788), .ZN(n783) );
  NR2D0 U50 ( .A1(port_dest[27]), .A2(n780), .ZN(n777) );
  AOI21D0 U51 ( .A1(n789), .A2(n790), .B(n734), .ZN(n780) );
  AN2D0 U52 ( .A1(n789), .A2(n791), .Z(n734) );
  OAI21D0 U53 ( .A1(n790), .A2(n792), .B(n793), .ZN(n791) );
  CKND0 U54 ( .I(n794), .ZN(n790) );
  MUX2ND0 U55 ( .I0(n360), .I1(n795), .S(n7), .ZN(n776) );
  MUX2ND0 U56 ( .I0(n361), .I1(n18), .S(n8), .ZN(n775) );
  CKND0 U57 ( .I(n796), .ZN(n18) );
  CKND0 U58 ( .I(n797), .ZN(n361) );
  MUX2ND0 U59 ( .I0(n798), .I1(n799), .S(n6), .ZN(N1616) );
  MUX3ND0 U60 ( .I0(n796), .I1(n797), .I2(n800), .S0(n8), .S1(n801), .ZN(N1615) );
  MUX2ND0 U61 ( .I0(n802), .I1(n358), .S(n7), .ZN(n800) );
  CKND0 U62 ( .I(n773), .ZN(n358) );
  INR2D0 U63 ( .A1(n803), .B1(n804), .ZN(n773) );
  MUX2ND0 U64 ( .I0(n805), .I1(\dst[5][1] ), .S(n806), .ZN(n803) );
  OAI22D0 U65 ( .A1(n807), .A2(n808), .B1(port_dest[11]), .B2(n809), .ZN(n805)
         );
  INR2D0 U66 ( .A1(n810), .B1(n811), .ZN(n809) );
  MUX2ND0 U67 ( .I0(n812), .I1(\dst[7][1] ), .S(n813), .ZN(n797) );
  IND2D0 U68 ( .A1(n814), .B1(n815), .ZN(n812) );
  OAI21D0 U69 ( .A1(n816), .A2(n817), .B(n818), .ZN(n815) );
  OAI22D0 U70 ( .A1(\dst[6][1] ), .A2(n819), .B1(n820), .B2(n821), .ZN(n796)
         );
  MUX2ND0 U71 ( .I0(n822), .I1(n823), .S(n824), .ZN(n821) );
  NR2D0 U72 ( .A1(n825), .A2(n826), .ZN(n823) );
  IAO21D0 U73 ( .A1(n827), .A2(n828), .B(n829), .ZN(n826) );
  MUX2ND0 U74 ( .I0(n799), .I1(n798), .S(n6), .ZN(N1614) );
  CKND0 U75 ( .I(n801), .ZN(n6) );
  XNR2D0 U76 ( .A1(n830), .A2(n20), .ZN(n801) );
  MUX2ND0 U77 ( .I0(n795), .I1(n360), .S(n7), .ZN(n830) );
  OAI21D0 U78 ( .A1(n831), .A2(n832), .B(n833), .ZN(n360) );
  MUX2ND0 U79 ( .I0(n834), .I1(\dst[5][2] ), .S(n806), .ZN(n833) );
  MUX2ND0 U80 ( .I0(n388), .I1(n386), .S(n8), .ZN(n798) );
  MUX4ND0 U81 ( .I0(n835), .I1(n836), .I2(n837), .I3(n838), .S0(n839), .S1(n19), .ZN(n8) );
  OA32D0 U82 ( .A1(n840), .A2(n841), .A3(n820), .B1(\dst[6][2] ), .B2(n819), 
        .Z(n19) );
  AOI31D0 U83 ( .A1(n842), .A2(n843), .A3(n844), .B(port_dest[7]), .ZN(n840)
         );
  OA22D0 U84 ( .A1(n845), .A2(n820), .B1(\dst[6][1] ), .B2(n819), .Z(n839) );
  MUX2D0 U85 ( .I0(n846), .I1(port_dest[5]), .S(port_dest[7]), .Z(n845) );
  OAI21D0 U86 ( .A1(n847), .A2(n829), .B(n843), .ZN(n846) );
  NR2D0 U87 ( .A1(n828), .A2(n827), .ZN(n847) );
  AN3D0 U88 ( .A1(n848), .A2(n849), .A3(n756), .Z(n838) );
  AN3D0 U89 ( .A1(n850), .A2(n851), .A3(n755), .Z(n837) );
  INR3D0 U90 ( .A1(n750), .B1(n751), .B2(n852), .ZN(n836) );
  NR3D0 U91 ( .A1(n853), .A2(n753), .A3(n854), .ZN(n835) );
  AO21D0 U92 ( .A1(\dst[7][0] ), .A2(n813), .B(n855), .Z(n386) );
  MUX2ND0 U93 ( .I0(n856), .I1(n857), .S(n818), .ZN(n855) );
  NR2D0 U94 ( .A1(n858), .A2(n859), .ZN(n857) );
  IINR4D0 U95 ( .A1(n860), .A2(n861), .B1(n816), .B2(n862), .ZN(n858) );
  IINR4D0 U96 ( .A1(n863), .A2(n864), .B1(n862), .B2(n859), .ZN(n813) );
  AN3D0 U97 ( .A1(n816), .A2(n865), .A3(n866), .Z(n859) );
  AOI221D0 U98 ( .A1(n867), .A2(n868), .B1(n869), .B2(n870), .C(n820), .ZN(
        n866) );
  NR2D0 U99 ( .A1(n868), .A2(n867), .ZN(n820) );
  IINR4D0 U100 ( .A1(n871), .A2(n872), .B1(n873), .B2(n874), .ZN(n816) );
  INR3D0 U101 ( .A1(n872), .B1(n873), .B2(n871), .ZN(n862) );
  OAI21D0 U102 ( .A1(port_dest[7]), .A2(n875), .B(n876), .ZN(n871) );
  AOI211D0 U103 ( .A1(n867), .A2(n868), .B(n817), .C(n877), .ZN(n864) );
  OAI21D0 U104 ( .A1(n872), .A2(n873), .B(n861), .ZN(n817) );
  OAI211D0 U105 ( .A1(port_dest[7]), .A2(n829), .B(n828), .C(n878), .ZN(n861)
         );
  OAI21D0 U106 ( .A1(n879), .A2(n880), .B(n878), .ZN(n873) );
  CKND0 U107 ( .I(n877), .ZN(n878) );
  CKND2D0 U108 ( .A1(n881), .A2(n860), .ZN(n877) );
  CKND2D0 U109 ( .A1(n882), .A2(port_dest[7]), .ZN(n860) );
  OAI21D0 U110 ( .A1(port_dest[7]), .A2(n882), .B(n883), .ZN(n881) );
  NR2D0 U111 ( .A1(port_dest[7]), .A2(n829), .ZN(n879) );
  OAI31D0 U112 ( .A1(n829), .A2(port_dest[7]), .A3(n828), .B(n827), .ZN(n872)
         );
  OR2D0 U113 ( .A1(n884), .A2(n885), .Z(n868) );
  NR2D0 U114 ( .A1(port_dest[3]), .A2(n874), .ZN(n863) );
  AN2D0 U115 ( .A1(n885), .A2(n884), .Z(n874) );
  CKND2D0 U116 ( .A1(n886), .A2(n824), .ZN(n884) );
  MUX3D0 U117 ( .I0(n887), .I1(port_dest[4]), .I2(\dst[6][0] ), .S0(
        port_dest[7]), .S1(n888), .Z(n388) );
  CKND0 U118 ( .I(n819), .ZN(n888) );
  ND4D0 U119 ( .A1(n843), .A2(n824), .A3(n842), .A4(n889), .ZN(n819) );
  AOI211D0 U120 ( .A1(n865), .A2(n890), .B(n875), .C(n891), .ZN(n889) );
  CKND0 U121 ( .I(n844), .ZN(n891) );
  CKND2D0 U122 ( .A1(n885), .A2(n886), .ZN(n844) );
  CKND2D0 U123 ( .A1(n869), .A2(n870), .ZN(n890) );
  INR4D0 U124 ( .A1(n842), .B1(n882), .B2(n825), .B3(n892), .ZN(n887) );
  NR2D0 U125 ( .A1(n829), .A2(n880), .ZN(n892) );
  CKND0 U126 ( .I(n843), .ZN(n825) );
  IND3D0 U127 ( .A1(n885), .B1(n886), .B2(n867), .ZN(n843) );
  NR2D0 U128 ( .A1(n870), .A2(n869), .ZN(n867) );
  NR2D0 U129 ( .A1(n810), .A2(port_dest[11]), .ZN(n869) );
  NR2D0 U130 ( .A1(n875), .A2(n876), .ZN(n886) );
  CKND0 U131 ( .I(n893), .ZN(n875) );
  AOI21D0 U132 ( .A1(n894), .A2(n834), .B(n895), .ZN(n885) );
  CKND2D0 U133 ( .A1(n876), .A2(n893), .ZN(n842) );
  NR3D0 U134 ( .A1(n827), .A2(n828), .A3(n829), .ZN(n893) );
  OR2D0 U135 ( .A1(n883), .A2(n882), .Z(n829) );
  NR2D0 U136 ( .A1(n896), .A2(n831), .ZN(n882) );
  NR2D0 U137 ( .A1(n897), .A2(n898), .ZN(n883) );
  CKND0 U138 ( .I(n880), .ZN(n828) );
  CKND2D0 U139 ( .A1(n899), .A2(n807), .ZN(n880) );
  IAO21D0 U140 ( .A1(n899), .A2(n807), .B(n808), .ZN(n827) );
  NR2D0 U141 ( .A1(n894), .A2(n834), .ZN(n876) );
  NR2D0 U142 ( .A1(n900), .A2(port_dest[11]), .ZN(n834) );
  MUX2ND0 U143 ( .I0(n901), .I1(n359), .S(n7), .ZN(n799) );
  AN3D0 U144 ( .A1(n848), .A2(n850), .A3(n902), .Z(n7) );
  AOI33D0 U145 ( .A1(n903), .A2(n852), .A3(n750), .B1(n904), .B2(n854), .B3(
        n752), .ZN(n902) );
  CKND0 U146 ( .I(n853), .ZN(n752) );
  OAI22D0 U147 ( .A1(\dst[2][2] ), .A2(n905), .B1(n376), .B2(n362), .ZN(n853)
         );
  OAI22D0 U148 ( .A1(n46), .A2(n277), .B1(\dst[4][1] ), .B2(n906), .ZN(n854)
         );
  CKND0 U149 ( .I(n907), .ZN(n906) );
  CKND0 U150 ( .I(n908), .ZN(n46) );
  CKND0 U151 ( .I(n753), .ZN(n904) );
  NR2D0 U152 ( .A1(n17), .A2(n20), .ZN(n753) );
  AOI32D0 U153 ( .A1(\dst[2][1] ), .A2(n909), .A3(n910), .B1(n911), .B2(n376), 
        .ZN(n750) );
  AO22D0 U154 ( .A1(n907), .A2(\dst[4][1] ), .B1(n908), .B2(n277), .Z(n852) );
  CKND0 U155 ( .I(n751), .ZN(n903) );
  NR2D0 U156 ( .A1(n912), .A2(n20), .ZN(n751) );
  ND3D0 U157 ( .A1(n755), .A2(n851), .A3(n913), .ZN(n850) );
  OAI32D0 U158 ( .A1(n914), .A2(\dst[4][1] ), .A3(n375), .B1(n277), .B2(n908), 
        .ZN(n913) );
  CKND0 U159 ( .I(\dst[4][2] ), .ZN(n914) );
  CKND2D0 U160 ( .A1(n851), .A2(n915), .ZN(n755) );
  OAI22D0 U161 ( .A1(n909), .A2(n905), .B1(n376), .B2(n911), .ZN(n915) );
  CKND2D0 U162 ( .A1(n20), .A2(n912), .ZN(n851) );
  CKND0 U163 ( .I(n17), .ZN(n912) );
  ND4D0 U164 ( .A1(n802), .A2(n795), .A3(n756), .A4(n849), .ZN(n848) );
  ND4D0 U165 ( .A1(n11), .A2(n849), .A3(n376), .A4(n905), .ZN(n756) );
  OR2D0 U166 ( .A1(\dst[2][1] ), .A2(n41), .Z(n905) );
  CKND0 U167 ( .I(n910), .ZN(n41) );
  OAI221D0 U168 ( .A1(n916), .A2(n917), .B1(n918), .B2(n919), .C(n920), .ZN(
        n376) );
  CKND2D0 U169 ( .A1(n17), .A2(n20), .ZN(n849) );
  ND3D0 U170 ( .A1(n921), .A2(n922), .A3(n923), .ZN(n20) );
  MAOI22D0 U171 ( .A1(\dst[0][2] ), .A2(n924), .B1(port_dest[31]), .B2(n925), 
        .ZN(n923) );
  OAI211D0 U172 ( .A1(n926), .A2(n927), .B(n921), .C(n928), .ZN(n17) );
  AOI21D0 U173 ( .A1(\dst[0][1] ), .A2(n924), .B(n929), .ZN(n928) );
  MUX2D0 U174 ( .I0(n717), .I1(port_dest[29]), .S(port_dest[31]), .Z(n929) );
  CKND0 U175 ( .I(n714), .ZN(n924) );
  CKND2D0 U176 ( .A1(n787), .A2(n714), .ZN(n921) );
  ND4D0 U177 ( .A1(n925), .A2(n930), .A3(n931), .A4(n927), .ZN(n714) );
  NR2D0 U178 ( .A1(n782), .A2(n717), .ZN(n931) );
  INR3D0 U179 ( .A1(n932), .B1(n933), .B2(n934), .ZN(n717) );
  CKND0 U180 ( .I(n935), .ZN(n782) );
  IAO21D0 U181 ( .A1(n936), .A2(n720), .B(n716), .ZN(n925) );
  INR3D0 U182 ( .A1(n936), .B1(n788), .B2(n720), .ZN(n716) );
  INR2D0 U183 ( .A1(n721), .B1(n937), .ZN(n936) );
  MUX2ND0 U184 ( .I0(n911), .I1(n909), .S(n910), .ZN(n11) );
  NR4D0 U185 ( .A1(n938), .A2(n748), .A3(n939), .A4(n940), .ZN(n910) );
  OA211D0 U186 ( .A1(n941), .A2(n942), .B(n943), .C(n916), .Z(n748) );
  NR3D0 U187 ( .A1(n792), .A2(n779), .A3(n940), .ZN(n942) );
  CKND0 U188 ( .I(\dst[2][2] ), .ZN(n909) );
  CKND0 U189 ( .I(n362), .ZN(n911) );
  IND2D0 U190 ( .A1(n944), .B1(n938), .ZN(n362) );
  NR2D0 U191 ( .A1(n908), .A2(n907), .ZN(n795) );
  NR2D0 U192 ( .A1(n375), .A2(\dst[4][2] ), .ZN(n907) );
  NR2D0 U193 ( .A1(n945), .A2(n946), .ZN(n908) );
  CKND0 U194 ( .I(n774), .ZN(n802) );
  OAI21D0 U195 ( .A1(\dst[4][1] ), .A2(n375), .B(n277), .ZN(n774) );
  OAI22D0 U196 ( .A1(n947), .A2(n948), .B1(n949), .B2(n950), .ZN(n277) );
  AOI211D0 U197 ( .A1(n951), .A2(n952), .B(n953), .C(n954), .ZN(n949) );
  OAI21D0 U198 ( .A1(n831), .A2(n955), .B(n956), .ZN(n359) );
  MUX2ND0 U199 ( .I0(n957), .I1(\dst[5][0] ), .S(n806), .ZN(n956) );
  NR4D0 U200 ( .A1(n958), .A2(n807), .A3(n811), .A4(n959), .ZN(n806) );
  CKND2D0 U201 ( .A1(n898), .A2(n897), .ZN(n807) );
  CKND0 U202 ( .I(n960), .ZN(n898) );
  IND3D0 U203 ( .A1(n865), .B1(n895), .B2(n808), .ZN(n958) );
  INR2D0 U204 ( .A1(n961), .B1(n758), .ZN(n865) );
  OAI21D0 U205 ( .A1(n962), .A2(n963), .B(n964), .ZN(n961) );
  NR3D0 U206 ( .A1(n959), .A2(n811), .A3(n960), .ZN(n957) );
  CKND2D0 U207 ( .A1(n896), .A2(n831), .ZN(n960) );
  AN3D0 U208 ( .A1(n897), .A2(n896), .A3(n899), .Z(n811) );
  CKND0 U209 ( .I(n965), .ZN(n899) );
  OAI22D0 U210 ( .A1(n900), .A2(n894), .B1(n810), .B2(n870), .ZN(n959) );
  OR2D0 U211 ( .A1(n964), .A2(n962), .Z(n870) );
  NR2D0 U212 ( .A1(n966), .A2(n967), .ZN(n962) );
  IND3D0 U213 ( .A1(n900), .B1(n895), .B2(n894), .ZN(n810) );
  CKND2D0 U214 ( .A1(n967), .A2(n966), .ZN(n895) );
  CKND2D0 U215 ( .A1(n946), .A2(n951), .ZN(n966) );
  CKND0 U216 ( .I(n968), .ZN(n951) );
  IND2D0 U217 ( .A1(n946), .B1(n968), .ZN(n894) );
  ND4D0 U218 ( .A1(n808), .A2(n965), .A3(n897), .A4(n896), .ZN(n900) );
  CKND2D0 U219 ( .A1(n969), .A2(port_dest[15]), .ZN(n896) );
  OAI21D0 U220 ( .A1(port_dest[15]), .A2(n969), .B(n970), .ZN(n897) );
  CKND2D0 U221 ( .A1(n953), .A2(n950), .ZN(n965) );
  OAI21D0 U222 ( .A1(n953), .A2(n950), .B(n954), .ZN(n808) );
  OA21D0 U223 ( .A1(\dst[4][0] ), .A2(n375), .B(n1), .Z(n901) );
  MUX2D0 U224 ( .I0(n971), .I1(port_dest[12]), .S(port_dest[15]), .Z(n1) );
  AOI211D0 U225 ( .A1(n953), .A2(n972), .B(n969), .C(n973), .ZN(n971) );
  CKND0 U226 ( .I(n974), .ZN(n973) );
  ND4D0 U227 ( .A1(n946), .A2(n975), .A3(n974), .A4(n952), .ZN(n375) );
  OAI211D0 U228 ( .A1(n968), .A2(n976), .B(n977), .C(n972), .ZN(n974) );
  CKND0 U229 ( .I(n954), .ZN(n977) );
  NR2D0 U230 ( .A1(n967), .A2(n964), .ZN(n976) );
  OR2D0 U231 ( .A1(n766), .A2(n978), .Z(n964) );
  CKND0 U232 ( .I(n952), .ZN(n967) );
  CKND2D0 U233 ( .A1(n760), .A2(n979), .ZN(n952) );
  NR2D0 U234 ( .A1(n767), .A2(n761), .ZN(n968) );
  OR2D0 U235 ( .A1(n963), .A2(n758), .Z(n975) );
  OAI21D0 U236 ( .A1(n980), .A2(n920), .B(n939), .ZN(n758) );
  AOI221D0 U237 ( .A1(n792), .A2(n779), .B1(n788), .B2(n787), .C(n935), .ZN(
        n939) );
  ND4D0 U238 ( .A1(n981), .A2(n982), .A3(n983), .A4(n984), .ZN(n935) );
  AOI33D0 U239 ( .A1(port_dest[4]), .A2(n841), .A3(port_dest[5]), .B1(
        port_dest[28]), .B2(n985), .B3(port_dest[29]), .ZN(n984) );
  AOI33D0 U240 ( .A1(port_dest[24]), .A2(n778), .A3(port_dest[25]), .B1(
        port_dest[20]), .B2(n944), .B3(port_dest[21]), .ZN(n983) );
  AOI33D0 U241 ( .A1(port_dest[16]), .A2(n762), .A3(port_dest[17]), .B1(
        port_dest[12]), .B2(n945), .B3(port_dest[13]), .ZN(n982) );
  AOI33D0 U242 ( .A1(port_dest[8]), .A2(port_dest[10]), .A3(n804), .B1(
        port_dest[2]), .B2(port_dest[0]), .B3(n814), .ZN(n981) );
  NR2D0 U243 ( .A1(n779), .A2(n792), .ZN(n980) );
  CKND0 U244 ( .I(n986), .ZN(n792) );
  CKND0 U245 ( .I(n727), .ZN(n779) );
  INR2D0 U246 ( .A1(n766), .B1(n757), .ZN(n963) );
  CKND0 U247 ( .I(n978), .ZN(n757) );
  NR2D0 U248 ( .A1(n979), .A2(n760), .ZN(n978) );
  INR2D0 U249 ( .A1(n940), .B1(n987), .ZN(n760) );
  CKND2D0 U250 ( .A1(n761), .A2(n767), .ZN(n979) );
  CKND2D0 U251 ( .A1(n941), .A2(n938), .ZN(n767) );
  INR2D0 U252 ( .A1(n764), .B1(port_dest[19]), .ZN(n761) );
  AN4D0 U253 ( .A1(n988), .A2(n742), .A3(n743), .A4(n739), .Z(n764) );
  ND3D0 U254 ( .A1(n920), .A2(n727), .A3(n986), .ZN(n766) );
  NR2D0 U255 ( .A1(n788), .A2(n787), .ZN(n986) );
  NR2D0 U256 ( .A1(n989), .A2(n937), .ZN(n787) );
  ND4D0 U257 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n788) );
  AOI33D0 U258 ( .A1(n944), .A2(n994), .A3(port_dest[21]), .B1(n762), .B2(n995), .B3(port_dest[17]), .ZN(n993) );
  AOI33D0 U259 ( .A1(n985), .A2(n719), .A3(port_dest[29]), .B1(n778), .B2(n735), .B3(port_dest[25]), .ZN(n992) );
  AOI33D0 U260 ( .A1(n841), .A2(n996), .A3(port_dest[5]), .B1(n945), .B2(n997), 
        .B3(port_dest[13]), .ZN(n991) );
  AOI33D0 U261 ( .A1(port_dest[2]), .A2(n856), .A3(n814), .B1(port_dest[10]), 
        .B2(n955), .B3(n804), .ZN(n990) );
  CKND2D0 U262 ( .A1(n998), .A2(n794), .ZN(n727) );
  IND2D0 U263 ( .A1(n940), .B1(n987), .ZN(n920) );
  NR2D0 U264 ( .A1(n938), .A2(n941), .ZN(n987) );
  AOI21D0 U265 ( .A1(n730), .A2(n789), .B(n793), .ZN(n941) );
  IND2D0 U266 ( .A1(n917), .B1(n916), .ZN(n938) );
  NR2D0 U267 ( .A1(n999), .A2(n745), .ZN(n916) );
  NR2D0 U268 ( .A1(n794), .A2(n998), .ZN(n940) );
  AN3D0 U269 ( .A1(n793), .A2(n730), .A3(n789), .Z(n998) );
  NR4D0 U270 ( .A1(n784), .A2(n1000), .A3(n749), .A4(n785), .ZN(n789) );
  OR2D0 U271 ( .A1(n721), .A2(n1001), .Z(n793) );
  CKND2D0 U272 ( .A1(n937), .A2(n989), .ZN(n794) );
  CKND2D0 U273 ( .A1(n1001), .A2(n721), .ZN(n989) );
  ND4D0 U274 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n721) );
  AOI33D0 U275 ( .A1(n1006), .A2(n955), .A3(port_dest[10]), .B1(n1007), .B2(
        n856), .B3(port_dest[2]), .ZN(n1005) );
  AOI33D0 U276 ( .A1(n994), .A2(n919), .A3(n944), .B1(n995), .B2(n1008), .B3(
        n762), .ZN(n1004) );
  AOI33D0 U277 ( .A1(n719), .A2(n1009), .A3(n985), .B1(n735), .B2(n1010), .B3(
        n778), .ZN(n1003) );
  AOI33D0 U278 ( .A1(n996), .A2(n822), .A3(n841), .B1(n997), .B2(n948), .B3(
        n945), .ZN(n1002) );
  NR2D0 U279 ( .A1(n720), .A2(port_dest[31]), .ZN(n1001) );
  ND4D0 U280 ( .A1(n927), .A2(n934), .A3(n932), .A4(n1011), .ZN(n720) );
  AN4D0 U281 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .Z(n937) );
  AOI33D0 U282 ( .A1(port_dest[10]), .A2(n1006), .A3(port_dest[8]), .B1(
        port_dest[0]), .B2(n1007), .B3(port_dest[2]), .ZN(n1015) );
  AOI33D0 U283 ( .A1(n944), .A2(n919), .A3(port_dest[20]), .B1(n762), .B2(
        n1008), .B3(port_dest[16]), .ZN(n1014) );
  AN2D0 U284 ( .A1(port_dest[18]), .A2(port_dest[19]), .Z(n762) );
  INR2D0 U285 ( .A1(port_dest[22]), .B1(n918), .ZN(n944) );
  AOI33D0 U286 ( .A1(n985), .A2(n1009), .A3(port_dest[28]), .B1(n778), .B2(
        n1010), .B3(port_dest[24]), .ZN(n1013) );
  AN2D0 U287 ( .A1(port_dest[26]), .A2(port_dest[27]), .Z(n778) );
  CKND0 U288 ( .I(n922), .ZN(n985) );
  CKND2D0 U289 ( .A1(port_dest[31]), .A2(port_dest[30]), .ZN(n922) );
  AOI33D0 U290 ( .A1(n841), .A2(n822), .A3(port_dest[4]), .B1(n945), .B2(n948), 
        .B3(port_dest[12]), .ZN(n1012) );
  INR2D0 U291 ( .A1(port_dest[14]), .B1(n947), .ZN(n945) );
  AN2D0 U292 ( .A1(port_dest[6]), .A2(port_dest[7]), .Z(n841) );
  NR3D0 U293 ( .A1(n954), .A2(n953), .A3(n950), .ZN(n946) );
  CKND2D0 U294 ( .A1(n972), .A2(n947), .ZN(n950) );
  NR2D0 U295 ( .A1(n970), .A2(n969), .ZN(n972) );
  NR2D0 U296 ( .A1(n742), .A2(n737), .ZN(n969) );
  AOI21D0 U297 ( .A1(n737), .A2(n742), .B(n743), .ZN(n970) );
  NR2D0 U298 ( .A1(n1016), .A2(n739), .ZN(n953) );
  AOI21D0 U299 ( .A1(n739), .A2(n1016), .B(n988), .ZN(n954) );
  OAI21D0 U300 ( .A1(n745), .A2(n917), .B(n999), .ZN(n988) );
  AOI21D0 U301 ( .A1(n786), .A2(n731), .B(n726), .ZN(n999) );
  CKND0 U302 ( .I(n784), .ZN(n726) );
  AOI21D0 U303 ( .A1(n934), .A2(n930), .B(n927), .ZN(n784) );
  ND4D0 U304 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n927) );
  AOI33D0 U305 ( .A1(n1021), .A2(port_dest[12]), .A3(port_dest[13]), .B1(n1022), .B2(port_dest[20]), .B3(port_dest[21]), .ZN(n1020) );
  AOI33D0 U306 ( .A1(n1023), .A2(port_dest[4]), .A3(port_dest[5]), .B1(n1024), 
        .B2(port_dest[16]), .B3(port_dest[17]), .ZN(n1019) );
  AOI33D0 U307 ( .A1(n1025), .A2(port_dest[24]), .A3(port_dest[25]), .B1(n1026), .B2(port_dest[28]), .B3(port_dest[29]), .ZN(n1018) );
  AOI33D0 U308 ( .A1(port_dest[0]), .A2(n1027), .A3(n814), .B1(port_dest[8]), 
        .B2(n832), .B3(n804), .ZN(n1017) );
  AN3D0 U309 ( .A1(n742), .A2(n743), .A3(n737), .Z(n1016) );
  OAI211D0 U310 ( .A1(port_dest[23]), .A2(n747), .B(n733), .C(n749), .ZN(n743)
         );
  CKND2D0 U311 ( .A1(n747), .A2(port_dest[23]), .ZN(n742) );
  CKND2D0 U312 ( .A1(n745), .A2(n917), .ZN(n739) );
  CKND2D0 U313 ( .A1(n943), .A2(n918), .ZN(n917) );
  AOI21D0 U314 ( .A1(n733), .A2(n749), .B(n747), .ZN(n943) );
  NR2D0 U315 ( .A1(n1028), .A2(n730), .ZN(n747) );
  NR2D0 U316 ( .A1(n786), .A2(n731), .ZN(n745) );
  NR2D0 U317 ( .A1(n733), .A2(n749), .ZN(n731) );
  NR2D0 U318 ( .A1(n932), .A2(n722), .ZN(n749) );
  CKND2D0 U319 ( .A1(n1028), .A2(n730), .ZN(n733) );
  CKND0 U320 ( .I(n785), .ZN(n1028) );
  NR2D0 U321 ( .A1(n1011), .A2(n718), .ZN(n785) );
  CKND0 U322 ( .I(n1000), .ZN(n786) );
  NR2D0 U323 ( .A1(n934), .A2(n930), .ZN(n1000) );
  CKND0 U324 ( .I(n926), .ZN(n930) );
  CKND2D0 U325 ( .A1(n722), .A2(n932), .ZN(n926) );
  ND4D0 U326 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n932) );
  AOI33D0 U327 ( .A1(port_dest[12]), .A2(n948), .A3(n1021), .B1(n1006), .B2(
        n832), .B3(port_dest[8]), .ZN(n1032) );
  AOI33D0 U328 ( .A1(port_dest[20]), .A2(n919), .A3(n1022), .B1(n1007), .B2(
        n1027), .B3(port_dest[0]), .ZN(n1031) );
  AOI33D0 U329 ( .A1(port_dest[4]), .A2(n822), .A3(n1023), .B1(port_dest[16]), 
        .B2(n1008), .B3(n1024), .ZN(n1030) );
  AOI33D0 U330 ( .A1(port_dest[24]), .A2(n1010), .A3(n1025), .B1(port_dest[28]), .B2(n1009), .B3(n1026), .ZN(n1029) );
  NR2D0 U331 ( .A1(n933), .A2(port_dest[31]), .ZN(n722) );
  CKND0 U332 ( .I(n1011), .ZN(n933) );
  ND4D0 U333 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1011) );
  AOI33D0 U334 ( .A1(n997), .A2(n948), .A3(n1021), .B1(n832), .B2(n955), .B3(
        n1006), .ZN(n1036) );
  NR2D0 U335 ( .A1(n831), .A2(port_dest[9]), .ZN(n1006) );
  CKND0 U336 ( .I(port_dest[13]), .ZN(n948) );
  AOI33D0 U337 ( .A1(n994), .A2(n919), .A3(n1022), .B1(n856), .B2(n1027), .B3(
        n1007), .ZN(n1035) );
  NR2D0 U338 ( .A1(n818), .A2(port_dest[1]), .ZN(n1007) );
  CKND0 U339 ( .I(port_dest[21]), .ZN(n919) );
  AOI33D0 U340 ( .A1(n996), .A2(n822), .A3(n1023), .B1(n995), .B2(n1008), .B3(
        n1024), .ZN(n1034) );
  CKND0 U341 ( .I(port_dest[17]), .ZN(n1008) );
  CKND0 U342 ( .I(port_dest[5]), .ZN(n822) );
  AOI33D0 U343 ( .A1(n735), .A2(n1010), .A3(n1025), .B1(n719), .B2(n1009), 
        .B3(n1026), .ZN(n1033) );
  CKND0 U344 ( .I(port_dest[29]), .ZN(n1009) );
  CKND0 U345 ( .I(port_dest[25]), .ZN(n1010) );
  ND4D0 U346 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n934) );
  AOI33D0 U347 ( .A1(n1021), .A2(n997), .A3(port_dest[13]), .B1(n1022), .B2(
        n994), .B3(port_dest[21]), .ZN(n1040) );
  CKND0 U348 ( .I(port_dest[20]), .ZN(n994) );
  NR2D0 U349 ( .A1(n918), .A2(port_dest[22]), .ZN(n1022) );
  CKND0 U350 ( .I(port_dest[23]), .ZN(n918) );
  CKND0 U351 ( .I(port_dest[12]), .ZN(n997) );
  NR2D0 U352 ( .A1(n947), .A2(port_dest[14]), .ZN(n1021) );
  CKND0 U353 ( .I(port_dest[15]), .ZN(n947) );
  AOI33D0 U354 ( .A1(n1023), .A2(n996), .A3(port_dest[5]), .B1(n1024), .B2(
        n995), .B3(port_dest[17]), .ZN(n1039) );
  CKND0 U355 ( .I(port_dest[16]), .ZN(n995) );
  NR2D0 U356 ( .A1(n737), .A2(port_dest[18]), .ZN(n1024) );
  CKND0 U357 ( .I(port_dest[19]), .ZN(n737) );
  CKND0 U358 ( .I(port_dest[4]), .ZN(n996) );
  NR2D0 U359 ( .A1(n824), .A2(port_dest[6]), .ZN(n1023) );
  CKND0 U360 ( .I(port_dest[7]), .ZN(n824) );
  AOI33D0 U361 ( .A1(n1025), .A2(n735), .A3(port_dest[25]), .B1(n1026), .B2(
        n719), .B3(port_dest[29]), .ZN(n1038) );
  CKND0 U362 ( .I(port_dest[28]), .ZN(n719) );
  NR2D0 U363 ( .A1(n718), .A2(port_dest[30]), .ZN(n1026) );
  CKND0 U364 ( .I(port_dest[31]), .ZN(n718) );
  CKND0 U365 ( .I(port_dest[24]), .ZN(n735) );
  NR2D0 U366 ( .A1(n730), .A2(port_dest[26]), .ZN(n1025) );
  CKND0 U367 ( .I(port_dest[27]), .ZN(n730) );
  AOI33D0 U368 ( .A1(n856), .A2(n1027), .A3(n814), .B1(n832), .B2(n955), .B3(
        n804), .ZN(n1037) );
  INR2D0 U369 ( .A1(port_dest[9]), .B1(n831), .ZN(n804) );
  CKND0 U370 ( .I(port_dest[11]), .ZN(n831) );
  CKND0 U371 ( .I(port_dest[8]), .ZN(n955) );
  CKND0 U372 ( .I(port_dest[10]), .ZN(n832) );
  INR2D0 U373 ( .A1(port_dest[1]), .B1(n818), .ZN(n814) );
  CKND0 U374 ( .I(port_dest[3]), .ZN(n818) );
  CKND0 U375 ( .I(port_dest[2]), .ZN(n1027) );
  CKND0 U376 ( .I(port_dest[0]), .ZN(n856) );
endmodule


module crossbar_0 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_4 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND2 U1 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND2 U2 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND2 U3 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND2 U4 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND2 U5 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND2 U6 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND2 U7 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND2 U8 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND2 U9 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND2 U10 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND2 U11 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND2 U12 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND2 U13 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND2 U14 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND2 U15 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND2 U16 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND2 U17 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND2 U18 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND2 U19 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND2 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND2 U21 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  MUX2ND2 U22 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  MUX2ND2 U23 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  MUX2ND2 U24 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  MUX2ND2 U25 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  MUX2ND2 U26 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  MUX2ND2 U27 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  MUX2ND2 U28 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  MUX2ND2 U29 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  MUX2ND2 U30 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  MUX2ND2 U31 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  MUX2ND2 U32 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  MUX2ND2 U33 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  MUX2ND2 U34 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  MUX2ND2 U35 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  MUX2ND2 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  MUX2ND2 U37 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  MUX2ND2 U38 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  MUX2ND2 U39 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  MUX2ND2 U40 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U41 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U42 ( .I(in_lower[9]), .ZN(n82) );
  CKND0 U43 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U44 ( .I(in_lower[8]), .ZN(n84) );
  CKND0 U45 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U46 ( .I(in_lower[7]), .ZN(n86) );
  CKND0 U47 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U48 ( .I(in_lower[6]), .ZN(n88) );
  CKND0 U49 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U50 ( .I(in_lower[5]), .ZN(n90) );
  CKND0 U51 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U52 ( .I(in_lower[4]), .ZN(n92) );
  CKND0 U53 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U54 ( .I(in_lower[3]), .ZN(n94) );
  CKND0 U55 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U56 ( .I(in_lower[2]), .ZN(n96) );
  CKND0 U57 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U58 ( .I(in_lower[1]), .ZN(n98) );
  CKND0 U59 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U60 ( .I(in_lower[19]), .ZN(n100) );
  CKND0 U61 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U62 ( .I(in_lower[18]), .ZN(n102) );
  CKND0 U63 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U64 ( .I(in_lower[17]), .ZN(n104) );
  CKND0 U65 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U66 ( .I(in_lower[16]), .ZN(n106) );
  CKND0 U67 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U68 ( .I(in_lower[15]), .ZN(n108) );
  CKND0 U69 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U70 ( .I(in_lower[14]), .ZN(n110) );
  CKND0 U71 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U72 ( .I(in_lower[13]), .ZN(n112) );
  CKND0 U73 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U74 ( .I(in_lower[12]), .ZN(n114) );
  CKND0 U75 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U76 ( .I(in_lower[11]), .ZN(n116) );
  CKND0 U77 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U78 ( .I(in_lower[10]), .ZN(n118) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_1 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND2 U1 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND2 U2 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND2 U3 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND2 U4 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND2 U5 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND2 U6 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND2 U7 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND2 U8 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND2 U9 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND2 U10 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND2 U11 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND2 U12 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND2 U13 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND2 U14 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND2 U15 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND2 U16 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND2 U17 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND2 U18 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND2 U19 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND2 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND2 U21 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  MUX2ND2 U22 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  MUX2ND2 U23 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  MUX2ND2 U24 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  MUX2ND2 U25 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  MUX2ND2 U26 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  MUX2ND2 U27 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  MUX2ND2 U28 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  MUX2ND2 U29 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  MUX2ND2 U30 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  MUX2ND2 U31 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  MUX2ND2 U32 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  MUX2ND2 U33 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  MUX2ND2 U34 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  MUX2ND2 U35 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  MUX2ND2 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  MUX2ND2 U37 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  MUX2ND2 U38 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  MUX2ND2 U39 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  MUX2ND2 U40 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U41 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U42 ( .I(in_lower[9]), .ZN(n82) );
  CKND0 U43 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U44 ( .I(in_lower[8]), .ZN(n84) );
  CKND0 U45 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U46 ( .I(in_lower[7]), .ZN(n86) );
  CKND0 U47 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U48 ( .I(in_lower[6]), .ZN(n88) );
  CKND0 U49 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U50 ( .I(in_lower[5]), .ZN(n90) );
  CKND0 U51 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U52 ( .I(in_lower[4]), .ZN(n92) );
  CKND0 U53 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U54 ( .I(in_lower[3]), .ZN(n94) );
  CKND0 U55 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U56 ( .I(in_lower[2]), .ZN(n96) );
  CKND0 U57 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U58 ( .I(in_lower[1]), .ZN(n98) );
  CKND0 U59 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U60 ( .I(in_lower[19]), .ZN(n100) );
  CKND0 U61 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U62 ( .I(in_lower[18]), .ZN(n102) );
  CKND0 U63 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U64 ( .I(in_lower[17]), .ZN(n104) );
  CKND0 U65 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U66 ( .I(in_lower[16]), .ZN(n106) );
  CKND0 U67 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U68 ( .I(in_lower[15]), .ZN(n108) );
  CKND0 U69 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U70 ( .I(in_lower[14]), .ZN(n110) );
  CKND0 U71 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U72 ( .I(in_lower[13]), .ZN(n112) );
  CKND0 U73 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U74 ( .I(in_lower[12]), .ZN(n114) );
  CKND0 U75 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U76 ( .I(in_lower[11]), .ZN(n116) );
  CKND0 U77 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U78 ( .I(in_lower[10]), .ZN(n118) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_2 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND2 U1 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND2 U2 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND2 U3 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND2 U4 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND2 U5 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND2 U6 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND2 U7 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND2 U8 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND2 U9 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND2 U10 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND2 U11 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND2 U12 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND2 U13 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND2 U14 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND2 U15 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND2 U16 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND2 U17 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND2 U18 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND2 U19 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND2 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND2 U21 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  MUX2ND2 U22 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  MUX2ND2 U23 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  MUX2ND2 U24 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  MUX2ND2 U25 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  MUX2ND2 U26 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  MUX2ND2 U27 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  MUX2ND2 U28 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  MUX2ND2 U29 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  MUX2ND2 U30 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  MUX2ND2 U31 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  MUX2ND2 U32 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  MUX2ND2 U33 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  MUX2ND2 U34 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  MUX2ND2 U35 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  MUX2ND2 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  MUX2ND2 U37 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  MUX2ND2 U38 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  MUX2ND2 U39 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  MUX2ND2 U40 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U41 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U42 ( .I(in_lower[9]), .ZN(n82) );
  CKND0 U43 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U44 ( .I(in_lower[8]), .ZN(n84) );
  CKND0 U45 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U46 ( .I(in_lower[7]), .ZN(n86) );
  CKND0 U47 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U48 ( .I(in_lower[6]), .ZN(n88) );
  CKND0 U49 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U50 ( .I(in_lower[5]), .ZN(n90) );
  CKND0 U51 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U52 ( .I(in_lower[4]), .ZN(n92) );
  CKND0 U53 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U54 ( .I(in_lower[3]), .ZN(n94) );
  CKND0 U55 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U56 ( .I(in_lower[2]), .ZN(n96) );
  CKND0 U57 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U58 ( .I(in_lower[1]), .ZN(n98) );
  CKND0 U59 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U60 ( .I(in_lower[19]), .ZN(n100) );
  CKND0 U61 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U62 ( .I(in_lower[18]), .ZN(n102) );
  CKND0 U63 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U64 ( .I(in_lower[17]), .ZN(n104) );
  CKND0 U65 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U66 ( .I(in_lower[16]), .ZN(n106) );
  CKND0 U67 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U68 ( .I(in_lower[15]), .ZN(n108) );
  CKND0 U69 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U70 ( .I(in_lower[14]), .ZN(n110) );
  CKND0 U71 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U72 ( .I(in_lower[13]), .ZN(n112) );
  CKND0 U73 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U74 ( .I(in_lower[12]), .ZN(n114) );
  CKND0 U75 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U76 ( .I(in_lower[11]), .ZN(n116) );
  CKND0 U77 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U78 ( .I(in_lower[10]), .ZN(n118) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_3 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND2 U1 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND2 U2 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND2 U3 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND2 U4 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND2 U5 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND2 U6 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND2 U7 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND2 U8 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND2 U9 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND2 U10 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND2 U11 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND2 U12 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND2 U13 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND2 U14 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND2 U15 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND2 U16 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND2 U17 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND2 U18 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND2 U19 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND2 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND2 U21 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  MUX2ND2 U22 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  MUX2ND2 U23 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  MUX2ND2 U24 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  MUX2ND2 U25 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  MUX2ND2 U26 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  MUX2ND2 U27 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  MUX2ND2 U28 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  MUX2ND2 U29 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  MUX2ND2 U30 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  MUX2ND2 U31 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  MUX2ND2 U32 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  MUX2ND2 U33 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  MUX2ND2 U34 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  MUX2ND2 U35 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  MUX2ND2 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  MUX2ND2 U37 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  MUX2ND2 U38 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  MUX2ND2 U39 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  MUX2ND2 U40 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U41 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U42 ( .I(in_lower[9]), .ZN(n82) );
  CKND0 U43 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U44 ( .I(in_lower[8]), .ZN(n84) );
  CKND0 U45 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U46 ( .I(in_lower[7]), .ZN(n86) );
  CKND0 U47 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U48 ( .I(in_lower[6]), .ZN(n88) );
  CKND0 U49 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U50 ( .I(in_lower[5]), .ZN(n90) );
  CKND0 U51 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U52 ( .I(in_lower[4]), .ZN(n92) );
  CKND0 U53 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U54 ( .I(in_lower[3]), .ZN(n94) );
  CKND0 U55 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U56 ( .I(in_lower[2]), .ZN(n96) );
  CKND0 U57 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U58 ( .I(in_lower[1]), .ZN(n98) );
  CKND0 U59 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U60 ( .I(in_lower[19]), .ZN(n100) );
  CKND0 U61 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U62 ( .I(in_lower[18]), .ZN(n102) );
  CKND0 U63 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U64 ( .I(in_lower[17]), .ZN(n104) );
  CKND0 U65 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U66 ( .I(in_lower[16]), .ZN(n106) );
  CKND0 U67 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U68 ( .I(in_lower[15]), .ZN(n108) );
  CKND0 U69 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U70 ( .I(in_lower[14]), .ZN(n110) );
  CKND0 U71 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U72 ( .I(in_lower[13]), .ZN(n112) );
  CKND0 U73 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U74 ( .I(in_lower[12]), .ZN(n114) );
  CKND0 U75 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U76 ( .I(in_lower[11]), .ZN(n116) );
  CKND0 U77 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U78 ( .I(in_lower[10]), .ZN(n118) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_5 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_6 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_7 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_8 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_9 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_10 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_11 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_12 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_13 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_14 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_15 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_16 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_17 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_18 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module crossbar_19 ( in_upper, in_lower, in_control, out_upper, out_lower );
  input [19:0] in_upper;
  input [19:0] in_lower;
  output [19:0] out_upper;
  output [19:0] out_lower;
  input in_control;
  wire   n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  MUX2ND0 U1 ( .I0(n81), .I1(n82), .S(in_control), .ZN(out_upper[9]) );
  MUX2ND0 U2 ( .I0(n83), .I1(n84), .S(in_control), .ZN(out_upper[8]) );
  MUX2ND0 U3 ( .I0(n85), .I1(n86), .S(in_control), .ZN(out_upper[7]) );
  MUX2ND0 U4 ( .I0(n87), .I1(n88), .S(in_control), .ZN(out_upper[6]) );
  MUX2ND0 U5 ( .I0(n89), .I1(n90), .S(in_control), .ZN(out_upper[5]) );
  MUX2ND0 U6 ( .I0(n91), .I1(n92), .S(in_control), .ZN(out_upper[4]) );
  MUX2ND0 U7 ( .I0(n93), .I1(n94), .S(in_control), .ZN(out_upper[3]) );
  MUX2ND0 U8 ( .I0(n95), .I1(n96), .S(in_control), .ZN(out_upper[2]) );
  MUX2ND0 U9 ( .I0(n97), .I1(n98), .S(in_control), .ZN(out_upper[1]) );
  MUX2ND0 U10 ( .I0(n99), .I1(n100), .S(in_control), .ZN(out_upper[19]) );
  MUX2ND0 U11 ( .I0(n101), .I1(n102), .S(in_control), .ZN(out_upper[18]) );
  MUX2ND0 U12 ( .I0(n103), .I1(n104), .S(in_control), .ZN(out_upper[17]) );
  MUX2ND0 U13 ( .I0(n105), .I1(n106), .S(in_control), .ZN(out_upper[16]) );
  MUX2ND0 U14 ( .I0(n107), .I1(n108), .S(in_control), .ZN(out_upper[15]) );
  MUX2ND0 U15 ( .I0(n109), .I1(n110), .S(in_control), .ZN(out_upper[14]) );
  MUX2ND0 U16 ( .I0(n111), .I1(n112), .S(in_control), .ZN(out_upper[13]) );
  MUX2ND0 U17 ( .I0(n113), .I1(n114), .S(in_control), .ZN(out_upper[12]) );
  MUX2ND0 U18 ( .I0(n115), .I1(n116), .S(in_control), .ZN(out_upper[11]) );
  MUX2ND0 U19 ( .I0(n117), .I1(n118), .S(in_control), .ZN(out_upper[10]) );
  MUX2ND0 U20 ( .I0(n119), .I1(n120), .S(in_control), .ZN(out_upper[0]) );
  MUX2ND0 U21 ( .I0(n82), .I1(n81), .S(in_control), .ZN(out_lower[9]) );
  CKND0 U22 ( .I(in_upper[9]), .ZN(n81) );
  CKND0 U23 ( .I(in_lower[9]), .ZN(n82) );
  MUX2ND0 U24 ( .I0(n84), .I1(n83), .S(in_control), .ZN(out_lower[8]) );
  CKND0 U25 ( .I(in_upper[8]), .ZN(n83) );
  CKND0 U26 ( .I(in_lower[8]), .ZN(n84) );
  MUX2ND0 U27 ( .I0(n86), .I1(n85), .S(in_control), .ZN(out_lower[7]) );
  CKND0 U28 ( .I(in_upper[7]), .ZN(n85) );
  CKND0 U29 ( .I(in_lower[7]), .ZN(n86) );
  MUX2ND0 U30 ( .I0(n88), .I1(n87), .S(in_control), .ZN(out_lower[6]) );
  CKND0 U31 ( .I(in_upper[6]), .ZN(n87) );
  CKND0 U32 ( .I(in_lower[6]), .ZN(n88) );
  MUX2ND0 U33 ( .I0(n90), .I1(n89), .S(in_control), .ZN(out_lower[5]) );
  CKND0 U34 ( .I(in_upper[5]), .ZN(n89) );
  CKND0 U35 ( .I(in_lower[5]), .ZN(n90) );
  MUX2ND0 U36 ( .I0(n92), .I1(n91), .S(in_control), .ZN(out_lower[4]) );
  CKND0 U37 ( .I(in_upper[4]), .ZN(n91) );
  CKND0 U38 ( .I(in_lower[4]), .ZN(n92) );
  MUX2ND0 U39 ( .I0(n94), .I1(n93), .S(in_control), .ZN(out_lower[3]) );
  CKND0 U40 ( .I(in_upper[3]), .ZN(n93) );
  CKND0 U41 ( .I(in_lower[3]), .ZN(n94) );
  MUX2ND0 U42 ( .I0(n96), .I1(n95), .S(in_control), .ZN(out_lower[2]) );
  CKND0 U43 ( .I(in_upper[2]), .ZN(n95) );
  CKND0 U44 ( .I(in_lower[2]), .ZN(n96) );
  MUX2ND0 U45 ( .I0(n98), .I1(n97), .S(in_control), .ZN(out_lower[1]) );
  CKND0 U46 ( .I(in_upper[1]), .ZN(n97) );
  CKND0 U47 ( .I(in_lower[1]), .ZN(n98) );
  MUX2ND0 U48 ( .I0(n100), .I1(n99), .S(in_control), .ZN(out_lower[19]) );
  CKND0 U49 ( .I(in_upper[19]), .ZN(n99) );
  CKND0 U50 ( .I(in_lower[19]), .ZN(n100) );
  MUX2ND0 U51 ( .I0(n102), .I1(n101), .S(in_control), .ZN(out_lower[18]) );
  CKND0 U52 ( .I(in_upper[18]), .ZN(n101) );
  CKND0 U53 ( .I(in_lower[18]), .ZN(n102) );
  MUX2ND0 U54 ( .I0(n104), .I1(n103), .S(in_control), .ZN(out_lower[17]) );
  CKND0 U55 ( .I(in_upper[17]), .ZN(n103) );
  CKND0 U56 ( .I(in_lower[17]), .ZN(n104) );
  MUX2ND0 U57 ( .I0(n106), .I1(n105), .S(in_control), .ZN(out_lower[16]) );
  CKND0 U58 ( .I(in_upper[16]), .ZN(n105) );
  CKND0 U59 ( .I(in_lower[16]), .ZN(n106) );
  MUX2ND0 U60 ( .I0(n108), .I1(n107), .S(in_control), .ZN(out_lower[15]) );
  CKND0 U61 ( .I(in_upper[15]), .ZN(n107) );
  CKND0 U62 ( .I(in_lower[15]), .ZN(n108) );
  MUX2ND0 U63 ( .I0(n110), .I1(n109), .S(in_control), .ZN(out_lower[14]) );
  CKND0 U64 ( .I(in_upper[14]), .ZN(n109) );
  CKND0 U65 ( .I(in_lower[14]), .ZN(n110) );
  MUX2ND0 U66 ( .I0(n112), .I1(n111), .S(in_control), .ZN(out_lower[13]) );
  CKND0 U67 ( .I(in_upper[13]), .ZN(n111) );
  CKND0 U68 ( .I(in_lower[13]), .ZN(n112) );
  MUX2ND0 U69 ( .I0(n114), .I1(n113), .S(in_control), .ZN(out_lower[12]) );
  CKND0 U70 ( .I(in_upper[12]), .ZN(n113) );
  CKND0 U71 ( .I(in_lower[12]), .ZN(n114) );
  MUX2ND0 U72 ( .I0(n116), .I1(n115), .S(in_control), .ZN(out_lower[11]) );
  CKND0 U73 ( .I(in_upper[11]), .ZN(n115) );
  CKND0 U74 ( .I(in_lower[11]), .ZN(n116) );
  MUX2ND0 U75 ( .I0(n118), .I1(n117), .S(in_control), .ZN(out_lower[10]) );
  CKND0 U76 ( .I(in_upper[10]), .ZN(n117) );
  CKND0 U77 ( .I(in_lower[10]), .ZN(n118) );
  MUX2ND0 U78 ( .I0(n120), .I1(n119), .S(in_control), .ZN(out_lower[0]) );
  CKND0 U79 ( .I(in_upper[0]), .ZN(n119) );
  CKND0 U80 ( .I(in_lower[0]), .ZN(n120) );
endmodule


module benes ( in_input, in_control, port_en_n, out_output );
  input [127:0] in_input;
  input [19:0] in_control;
  input [7:0] port_en_n;
  output [159:0] out_output;
  wire   \in_upper_00[3] , \in_lower_00[3] , \in_upper_01[3] ,
         \in_lower_01[3] , in_upper_02_3, \in_lower_02[3] , \in_upper_03[3] ,
         n1;
  wire   [19:0] in_upper_10;
  wire   [19:0] in_upper_12;
  wire   [19:0] in_lower_10;
  wire   [19:0] in_lower_12;
  wire   [19:0] in_upper_11;
  wire   [19:0] in_upper_13;
  wire   [19:0] in_lower_11;
  wire   [19:0] in_lower_13;
  wire   [19:0] in_upper_20;
  wire   [19:0] in_upper_21;
  wire   [19:0] in_lower_20;
  wire   [19:0] in_lower_21;
  wire   [19:0] in_upper_22;
  wire   [19:0] in_upper_23;
  wire   [19:0] in_lower_22;
  wire   [19:0] in_lower_23;
  wire   [19:0] in_upper_30;
  wire   [19:0] in_upper_31;
  wire   [19:0] in_lower_30;
  wire   [19:0] in_lower_31;
  wire   [19:0] in_upper_32;
  wire   [19:0] in_upper_33;
  wire   [19:0] in_lower_32;
  wire   [19:0] in_lower_33;
  wire   [19:0] in_upper_40;
  wire   [19:0] in_upper_41;
  wire   [19:0] in_upper_42;
  wire   [19:0] in_upper_43;
  wire   [19:0] in_lower_40;
  wire   [19:0] in_lower_41;
  wire   [19:0] in_lower_42;
  wire   [19:0] in_lower_43;
  assign \in_upper_00[3]  = port_en_n[0];
  assign \in_lower_00[3]  = port_en_n[1];
  assign \in_upper_01[3]  = port_en_n[2];
  assign \in_lower_01[3]  = port_en_n[3];
  assign in_upper_02_3 = port_en_n[4];
  assign \in_lower_02[3]  = port_en_n[5];
  assign \in_upper_03[3]  = port_en_n[6];

  crossbar_0 u_00_crossbar ( .in_upper({in_input[127:112], \in_upper_00[3] , 
        \in_upper_00[3] , \in_upper_00[3] , \in_upper_00[3] }), .in_lower({
        in_input[111:96], \in_lower_00[3] , \in_lower_00[3] , \in_lower_00[3] , 
        n1}), .in_control(in_control[19]), .out_upper(in_upper_10), 
        .out_lower(in_upper_12) );
  crossbar_19 u_01_crossbar ( .in_upper({in_input[95:80], \in_upper_01[3] , 
        \in_upper_01[3] , n1, \in_upper_01[3] }), .in_lower({in_input[79:64], 
        \in_lower_01[3] , \in_lower_01[3] , n1, n1}), .in_control(
        in_control[18]), .out_upper(in_lower_10), .out_lower(in_lower_12) );
  crossbar_18 u_02_crossbar ( .in_upper({in_input[63:48], in_upper_02_3, n1, 
        in_upper_02_3, in_upper_02_3}), .in_lower({in_input[47:32], 
        \in_lower_02[3] , n1, \in_lower_02[3] , n1}), .in_control(
        in_control[17]), .out_upper(in_upper_11), .out_lower(in_upper_13) );
  crossbar_17 u_03_crossbar ( .in_upper({in_input[31:16], \in_upper_03[3] , n1, 
        n1, \in_upper_03[3] }), .in_lower({in_input[15:0], port_en_n[7], n1, 
        n1, n1}), .in_control(in_control[16]), .out_upper(in_lower_11), 
        .out_lower(in_lower_13) );
  crossbar_16 u_10_crossbar ( .in_upper(in_upper_10), .in_lower(in_lower_10), 
        .in_control(in_control[15]), .out_upper(in_upper_20), .out_lower(
        in_upper_21) );
  crossbar_15 u_11_crossbar ( .in_upper(in_upper_11), .in_lower(in_lower_11), 
        .in_control(in_control[14]), .out_upper(in_lower_20), .out_lower(
        in_lower_21) );
  crossbar_14 u_12_crossbar ( .in_upper(in_upper_12), .in_lower(in_lower_12), 
        .in_control(in_control[13]), .out_upper(in_upper_22), .out_lower(
        in_upper_23) );
  crossbar_13 u_13_crossbar ( .in_upper(in_upper_13), .in_lower(in_lower_13), 
        .in_control(in_control[12]), .out_upper(in_lower_22), .out_lower(
        in_lower_23) );
  crossbar_12 u_20_crossbar ( .in_upper(in_upper_20), .in_lower(in_lower_20), 
        .in_control(in_control[11]), .out_upper(in_upper_30), .out_lower(
        in_upper_31) );
  crossbar_11 u_21_crossbar ( .in_upper(in_upper_21), .in_lower(in_lower_21), 
        .in_control(in_control[10]), .out_upper(in_lower_30), .out_lower(
        in_lower_31) );
  crossbar_10 u_22_crossbar ( .in_upper(in_upper_22), .in_lower(in_lower_22), 
        .in_control(in_control[9]), .out_upper(in_upper_32), .out_lower(
        in_upper_33) );
  crossbar_9 u_23_crossbar ( .in_upper(in_upper_23), .in_lower(in_lower_23), 
        .in_control(in_control[8]), .out_upper(in_lower_32), .out_lower(
        in_lower_33) );
  crossbar_8 u_30_crossbar ( .in_upper(in_upper_30), .in_lower(in_lower_30), 
        .in_control(in_control[7]), .out_upper(in_upper_40), .out_lower(
        in_upper_41) );
  crossbar_7 u_31_crossbar ( .in_upper(in_upper_31), .in_lower(in_lower_31), 
        .in_control(in_control[6]), .out_upper(in_upper_42), .out_lower(
        in_upper_43) );
  crossbar_6 u_32_crossbar ( .in_upper(in_upper_32), .in_lower(in_lower_32), 
        .in_control(in_control[5]), .out_upper(in_lower_40), .out_lower(
        in_lower_41) );
  crossbar_5 u_33_crossbar ( .in_upper(in_upper_33), .in_lower(in_lower_33), 
        .in_control(in_control[4]), .out_upper(in_lower_42), .out_lower(
        in_lower_43) );
  crossbar_4 u_40_crossbar ( .in_upper(in_upper_40), .in_lower(in_lower_40), 
        .in_control(in_control[3]), .out_upper(out_output[159:140]), 
        .out_lower(out_output[139:120]) );
  crossbar_3 u_41_crossbar ( .in_upper(in_upper_41), .in_lower(in_lower_41), 
        .in_control(in_control[2]), .out_upper(out_output[119:100]), 
        .out_lower(out_output[99:80]) );
  crossbar_2 u_42_crossbar ( .in_upper(in_upper_42), .in_lower(in_lower_42), 
        .in_control(in_control[1]), .out_upper(out_output[79:60]), .out_lower(
        out_output[59:40]) );
  crossbar_1 u_43_crossbar ( .in_upper(in_upper_43), .in_lower(in_lower_43), 
        .in_control(in_control[0]), .out_upper(out_output[39:20]), .out_lower(
        out_output[19:0]) );
  TIEH U3 ( .Z(n1) );
endmodule


module router ( clk, rst, fwd_routing_engine_port_dest, fwd_benes_out_output, 
        fwd_routing_engine_done );
  input [31:0] fwd_routing_engine_port_dest;
  output [159:0] fwd_benes_out_output;
  input clk, rst;
  output fwd_routing_engine_done;
  wire   n7;
  wire   [19:0] fwd_routing_engine_control;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  routing_engine_CLOCKED u_fwd_routing_engine ( .port_dest(
        fwd_routing_engine_port_dest), .clk(clk), .rst(rst), .control({
        SYNOPSYS_UNCONNECTED__0, fwd_routing_engine_control[18:16], 
        SYNOPSYS_UNCONNECTED__1, fwd_routing_engine_control[14], 
        SYNOPSYS_UNCONNECTED__2, fwd_routing_engine_control[12:0]}) );
  benes u_fwd_benes ( .in_input({n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, n7, n7, n7, n7, n7, n7, n7, n7}), .in_control({n7, 
        fwd_routing_engine_control[18:16], n7, fwd_routing_engine_control[14], 
        n7, fwd_routing_engine_control[12:0]}), .port_en_n({
        fwd_routing_engine_port_dest[3], fwd_routing_engine_port_dest[7], 
        fwd_routing_engine_port_dest[11], fwd_routing_engine_port_dest[15], 
        fwd_routing_engine_port_dest[19], fwd_routing_engine_port_dest[23], 
        fwd_routing_engine_port_dest[27], fwd_routing_engine_port_dest[31]}), 
        .out_output(fwd_benes_out_output) );
  TIEL U5 ( .ZN(n7) );
  TIEH U6 ( .Z(fwd_routing_engine_done) );
endmodule

