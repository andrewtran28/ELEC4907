module fma_mult_tree
  (
   input logic [9:0] mantissa_a,
   input logic [9:0] mantissa_b,
   input logic       sign_a,
   input logic       sign_b,

   output logic [19:0] mantissa_ab,
   output logic        sign_ab
   );

   logic [19:0]      x;
   logic [9:0]       y;
   logic [19:0]      pp0;
   logic [17:0]      pp1;
   logic [15:0]      pp2;
   logic [13:0]      pp3;
   logic [11:0]      pp4;
   logic [9:0]       pp5;
   logic [19:0]      int1, int2, p, g, c;
   logic [4:0][19:0] gp;
   logic [3:0][19:0] pp;
   logic [62:0][1:0] s;

   assign sign_ab = sign_a ^ sign_b;
   
   always_comb begin
      x = {10'h0, mantissa_a};
      y = mantissa_b;

      // Partial products
      pp0 = ((({20{y[0]^1'b0}} & x) | ({20{y[1]&~y[0]}} & {x[18:0],1'b0})) ^ {20{y[1]}}) + y[1];
      pp1 = ((({18{y[2]^y[1]}} & x[17:0]) | ({18{(~y[3]&y[2]&y[1])|(y[3]&~y[2]&~y[1])}} & {x[16:0],1'b0})) ^ {18{y[3]}}) + y[3];
      pp2 = ((({16{y[4]^y[3]}} & x[15:0]) | ({16{(~y[5]&y[4]&y[3])|(y[5]&~y[4]&~y[3])}} & {x[14:0],1'b0})) ^ {16{y[5]}}) + y[5];
      pp3 = ((({14{y[6]^y[5]}} & x[13:0]) | ({14{(~y[7]&y[6]&y[5])|(y[7]&~y[6]&~y[5])}} & {x[12:0],1'b0})) ^ {14{y[7]}}) + y[7];
      pp4 = ((({12{y[8]^y[7]}} & x[11:0]) | ({12{(~y[9]&y[8]&y[7])|(y[9]&~y[8]&~y[7])}} & {x[10:0],1'b0})) ^ {12{y[9]}}) + y[9];
      pp5 = {10{y[9]}} & x[9:0];

      // Wallace tree reduction layer 1
      s[0]  = pp0[2]+pp1[0];
      s[1]  = pp0[3]+pp1[1];
      s[2]  = pp0[4]+pp1[2]+pp2[0];
      s[3]  = pp0[5]+pp1[3]+pp2[1];
      s[4]  = pp0[6]+pp1[4]+pp2[2];
      s[5]  = pp0[7]+pp1[5]+pp2[3];
      s[6]  = pp0[8]+pp1[6]+pp2[4];
      s[7]  = pp3[2]+pp4[0];
      s[8]  = pp0[9]+pp1[7]+pp2[5];
      s[9]  = pp3[3]+pp4[1];
      s[10] = pp0[10]+pp1[8]+pp2[6];
      s[11] = pp3[4]+pp4[2]+pp5[0];
      s[12] = pp0[11]+pp1[9]+pp2[7];
      s[13] = pp3[5]+pp4[3]+pp5[1];
      s[14] = pp0[12]+pp1[10]+pp2[8];
      s[15] = pp3[6]+pp4[4]+pp5[2];
      s[16] = pp0[13]+pp1[11]+pp2[9];
      s[17] = pp3[7]+pp4[5]+pp5[3];
      s[18] = pp0[14]+pp1[12]+pp2[10];
      s[19] = pp3[8]+pp4[6]+pp5[4];
      s[20] = pp0[15]+pp1[13]+pp2[11];
      s[21] = pp3[9]+pp4[7]+pp5[5];
      s[22] = pp0[16]+pp1[14]+pp2[12];
      s[23] = pp3[10]+pp4[8]+pp5[6];
      s[24] = pp0[17]+pp1[15]+pp2[13];
      s[25] = pp3[11]+pp4[9]+pp5[7];
      s[26] = pp0[18]+pp1[16]+pp2[14];
      s[27] = pp3[12]+pp4[10]+pp5[8];
      s[28] = pp0[19]+pp1[17]+pp2[15];
      s[29] = pp3[13]+pp4[11]+pp5[9];

      // Wallace tree reduction layer 2
      s[30] = s[1][0]+s[0][1];
      s[31] = s[2][0]+s[1][1];
      s[32] = s[3][0]+s[2][1];
      s[33] = s[4][0]+s[3][1]+pp3[0];
      s[34] = s[5][0]+s[4][1]+pp3[1];
      s[35] = s[6][0]+s[7][0]+s[5][1];
      s[36] = s[8][0]+s[9][0]+s[6][1];
      s[37] = s[10][0]+s[11][0]+s[8][1];
      s[38] = s[12][0]+s[13][0]+s[10][1];
      s[39] = s[14][0]+s[15][0]+s[12][1];
      s[40] = s[16][0]+s[17][0]+s[14][1];
      s[41] = s[18][0]+s[19][0]+s[16][1];
      s[42] = s[20][0]+s[21][0]+s[18][1];
      s[43] = s[22][0]+s[23][0]+s[20][1];
      s[44] = s[24][0]+s[25][0]+s[22][1];
      s[45] = s[26][0]+s[27][0]+s[24][1];
      s[46] = s[28][0]+s[29][0]+s[26][1];

      // Wallace tree reduction layer 3
      s[47] = s[31][0]+s[30][1];
      s[48] = s[32][0]+s[31][1];
      s[49] = s[33][0]+s[32][1];
      s[50] = s[34][0]+s[33][1];
      s[51] = s[35][0]+s[34][1];
      s[52] = s[36][0]+s[35][1]+s[7][1];
      s[53] = s[37][0]+s[36][1]+s[9][1];
      s[54] = s[38][0]+s[37][1]+s[11][1];
      s[55] = s[39][0]+s[38][1]+s[13][1];
      s[56] = s[40][0]+s[39][1]+s[15][1];
      s[57] = s[41][0]+s[40][1]+s[17][1];
      s[58] = s[42][0]+s[41][1]+s[19][1];
      s[59] = s[43][0]+s[42][1]+s[21][1];
      s[60] = s[44][0]+s[43][1]+s[23][1];
      s[61] = s[45][0]+s[44][1]+s[25][1];
      s[62] = s[46][0]+s[45][1]+s[27][1];

      int1 = {s[62][0],s[61][0],s[60][0],s[59][0],s[58][0],s[57][0],s[56][0],s[55][0],s[54][0],s[53][0],s[52][0],s[51][0],s[50][0],s[49][0],s[48][0],s[47][0],s[30][0],s[0][0],pp0[1],pp0[0]};
      int2 = {s[61][1],s[60][1],s[59][1],s[58][1],s[57][1],s[56][1],s[55][1],s[54][1],s[53][1],s[52][1],s[51][1],s[50][1],s[49][1],s[48][1],s[47][1],1'b0    ,1'b0    ,1'b0   ,1'b0  ,1'b0  };

      // 20-bit Kogge-Stone Adder
      for (int i=0; i<20; i++) begin
         p[i] = int1[i]^int2[i];
         g[i] = int1[i]&int2[i];
      end

      pp[0][0] = p[0];
      gp[0][0] = g[0];
      for (int i=1; i<20; i++) begin
         pp[0][i] = p[i]&p[i-1];
         gp[0][i] = (p[i]&g[i-1])|g[i];
      end

      pp[1][0] = pp[0][0];
      pp[1][1] = pp[0][1];
      gp[1][0] = gp[0][0];
      gp[1][1] = gp[0][1];
      for (int i=2; i<20; i++) begin
         pp[1][i] = pp[0][i]&pp[0][i-2];
         gp[1][i] = (pp[0][i]&gp[0][i-2])|gp[0][i];
      end

      pp[2][0] = gp[1][0];
      pp[2][1] = gp[1][1];
      pp[2][2] = gp[1][2];
      pp[2][3] = gp[1][3];
      gp[2][0] = gp[1][0];
      gp[2][1] = gp[1][1];
      gp[2][2] = gp[1][2];
      gp[2][3] = gp[1][3];
      for (int i=4; i<20; i++) begin
         pp[2][i] = pp[1][i]&pp[1][i-4];
         gp[2][i] = (pp[1][i]&gp[1][i-4])|gp[1][i];
      end

      pp[3][0] = pp[2][0];
      pp[3][1] = pp[2][1];
      pp[3][2] = pp[2][2];
      pp[3][3] = pp[2][3];
      pp[3][4] = pp[2][4];
      pp[3][5] = pp[2][5];
      pp[3][6] = pp[2][6];
      pp[3][7] = pp[2][7];
      gp[3][0] = gp[2][0];
      gp[3][1] = gp[2][1];
      gp[3][2] = gp[2][2];
      gp[3][3] = gp[2][3];
      gp[3][4] = gp[2][4];
      gp[3][5] = gp[2][5];
      gp[3][6] = gp[2][6];
      gp[3][7] = gp[2][7];
      for (int i=8; i<20; i++) begin
         pp[3][i] = pp[2][i]&pp[2][i-8];
         gp[3][i] = (pp[2][i]&gp[2][i-8])|gp[2][i];
      end

      gp[4][0]  = gp[3][0];
      gp[4][1]  = gp[3][1];
      gp[4][2]  = gp[3][2];
      gp[4][3]  = gp[3][3];
      gp[4][4]  = gp[3][4];
      gp[4][5]  = gp[3][5];
      gp[4][6]  = gp[3][6];
      gp[4][7]  = gp[3][7];
      gp[4][8]  = gp[3][8];
      gp[4][9]  = gp[3][9];
      gp[4][10] = gp[3][10];
      gp[4][11] = gp[3][11];
      gp[4][12] = gp[3][12];
      gp[4][13] = gp[3][13];
      gp[4][14] = gp[3][14];
      gp[4][15] = gp[3][15];
      for (int i=16; i<20; i++) begin
         gp[4][i] = (pp[3][i]&gp[3][i-16])|gp[3][i];
      end

      mantissa_ab[0] = p[0];
      c[0]           = gp[4][0];
      for (int i=1; i<20; i++) begin
         mantissa_ab[i] = p[i]^c[i-1];
         c[i]           = gp[4][i];
      end
   end // always_comb

endmodule // fma_mult_tree