
module RamChip ( Address, Data, CS, WE, OE, clk, rst );
  input [6:0] Address;
  inout [47:0] Data;
  input CS, WE, OE, clk, rst;
  wire   \Mem[44][47] , \Mem[44][46] , \Mem[44][45] , \Mem[44][44] ,
         \Mem[44][43] , \Mem[44][42] , \Mem[44][41] , \Mem[44][40] ,
         \Mem[44][39] , \Mem[44][38] , \Mem[44][37] , \Mem[44][36] ,
         \Mem[44][35] , \Mem[44][34] , \Mem[44][33] , \Mem[44][32] ,
         \Mem[44][31] , \Mem[44][30] , \Mem[44][29] , \Mem[44][28] ,
         \Mem[44][27] , \Mem[44][26] , \Mem[44][25] , \Mem[44][24] ,
         \Mem[44][23] , \Mem[44][22] , \Mem[44][21] , \Mem[44][20] ,
         \Mem[44][19] , \Mem[44][18] , \Mem[44][17] , \Mem[44][16] ,
         \Mem[44][15] , \Mem[44][14] , \Mem[44][13] , \Mem[44][12] ,
         \Mem[44][11] , \Mem[44][10] , \Mem[44][9] , \Mem[44][8] ,
         \Mem[44][7] , \Mem[44][6] , \Mem[44][5] , \Mem[44][4] , \Mem[44][3] ,
         \Mem[44][2] , \Mem[44][1] , \Mem[44][0] , \Mem[45][47] ,
         \Mem[45][46] , \Mem[45][45] , \Mem[45][44] , \Mem[45][43] ,
         \Mem[45][42] , \Mem[45][41] , \Mem[45][40] , \Mem[45][39] ,
         \Mem[45][38] , \Mem[45][37] , \Mem[45][36] , \Mem[45][35] ,
         \Mem[45][34] , \Mem[45][33] , \Mem[45][32] , \Mem[45][31] ,
         \Mem[45][30] , \Mem[45][29] , \Mem[45][28] , \Mem[45][27] ,
         \Mem[45][26] , \Mem[45][25] , \Mem[45][24] , \Mem[45][23] ,
         \Mem[45][22] , \Mem[45][21] , \Mem[45][20] , \Mem[45][19] ,
         \Mem[45][18] , \Mem[45][17] , \Mem[45][16] , \Mem[45][15] ,
         \Mem[45][14] , \Mem[45][13] , \Mem[45][12] , \Mem[45][11] ,
         \Mem[45][10] , \Mem[45][9] , \Mem[45][8] , \Mem[45][7] , \Mem[45][6] ,
         \Mem[45][5] , \Mem[45][4] , \Mem[45][3] , \Mem[45][2] , \Mem[45][1] ,
         \Mem[45][0] , n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6460, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6477, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n15448, n15449, n15452, n15453,
         n15456, n15457, n15460, n15461, n15464, n15465, n15468, n15469,
         n15472, n15473, n15476, n15477, n15480, n15481, n15484, n15485,
         n15488, n15489, n15492, n15493, n15496, n15497, n15500, n15501,
         n15504, n15505, n15508, n15509, n15512, n15513, n15516, n15517,
         n15520, n15521, n15524, n15525, n15528, n15529, n15532, n15533,
         n15536, n15537, n15540, n15541, n15544, n15545, n15548, n15549,
         n15552, n15553, n15556, n15557, n15560, n15561, n15564, n15565,
         n15568, n15569, n15572, n15573, n15576, n15577, n15580, n15581,
         n15584, n15585, n15588, n15589, n15592, n15593, n15596, n15597,
         n15600, n15601, n15604, n15605, n15608, n15609, n15612, n15613,
         n15616, n15617, n15620, n15621, n15624, n15625, n15628, n15629,
         n15632, n15633, n15636, n15637, n15642, n17926, n17927, n17929,
         n17930, n17932, n17933, n17935, n17936, n17938, n17939, n17941,
         n17942, n17944, n17945, n17947, n17948, n17950, n17951, n17953,
         n17954, n17956, n17957, n17959, n17960, n17962, n17963, n17965,
         n17966, n17968, n17969, n17971, n17972, n17974, n17975, n17977,
         n17978, n17980, n17981, n17983, n17984, n17986, n17987, n17989,
         n17990, n17992, n17993, n17995, n17996, n17998, n17999, n18001,
         n18002, n18004, n18005, n18007, n18008, n18010, n18011, n18013,
         n18014, n18016, n18017, n18019, n18020, n18022, n18023, n18025,
         n18026, n18028, n18029, n18031, n18032, n18034, n18035, n18037,
         n18038, n18040, n18041, n18043, n18044, n18046, n18047, n18049,
         n18050, n18052, n18053, n18055, n18056, n18058, n18059, n18061,
         n18062, n18064, n18065, n18067, n18068, n24559, n24562, n24565,
         n24568, n24571, n24574, n24577, n24580, n24583, n24586, n24589,
         n24592, n24595, n24598, n24601, n24604, n24607, n24610, n24613,
         n24616, n24619, n24622, n24625, n24628, n24631, n24634, n24637,
         n24640, n24643, n24646, n24649, n24652, n24655, n24658, n24661,
         n24664, n24667, n24670, n24673, n24676, n24679, n24682, n24685,
         n24688, n24691, n24694, n24697, n24700, n24703, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227;
  tri   n15660;
  tri   n15662;
  tri   n15664;
  tri   n15666;
  tri   n15668;
  tri   n15670;
  tri   n15672;
  tri   n15674;
  tri   n15676;
  tri   n15678;
  tri   n15680;
  tri   n15682;
  tri   n15684;
  tri   n15686;
  tri   n15688;
  tri   n15690;
  tri   n15692;
  tri   n15694;
  tri   n15696;
  tri   n15698;
  tri   n15700;
  tri   n15702;
  tri   n15704;
  tri   n15706;
  tri   n15708;
  tri   n15710;
  tri   n15712;
  tri   n15714;
  tri   n15716;
  tri   n15718;
  tri   n15720;
  tri   n15722;
  tri   n15724;
  tri   n15726;
  tri   n15728;
  tri   n15730;
  tri   n15732;
  tri   n15734;
  tri   n15736;
  tri   n15738;
  tri   n15740;
  tri   n15742;
  tri   n15744;
  tri   n15746;
  tri   n15748;
  tri   n15750;
  tri   n15752;
  tri   n15754;
/*
  tran( n15660, Data[0]);
  tran( n15662, Data[1]);
  tran( n15664, Data[2]);
  tran( n15666, Data[3]);
  tran( n15668, Data[4]);
  tran( n15670, Data[5]);
  tran( n15672, Data[6]);
  tran( n15674, Data[7]);
  tran( n15676, Data[8]);
  tran( n15678, Data[9]);
  tran( n15680, Data[10]);
  tran( n15682, Data[11]);
  tran( n15684, Data[12]);
  tran( n15686, Data[13]);
  tran( n15688, Data[14]);
  tran( n15690, Data[15]);
  tran( n15692, Data[16]);
  tran( n15694, Data[17]);
  tran( n15696, Data[18]);
  tran( n15698, Data[19]);
  tran( n15700, Data[20]);
  tran( n15702, Data[21]);
  tran( n15704, Data[22]);
  tran( n15706, Data[23]);
  tran( n15708, Data[24]);
  tran( n15710, Data[25]);
  tran( n15712, Data[26]);
  tran( n15714, Data[27]);
  tran( n15716, Data[28]);
  tran( n15718, Data[29]);
  tran( n15720, Data[30]);
  tran( n15722, Data[31]);
  tran( n15724, Data[32]);
  tran( n15726, Data[33]);
  tran( n15728, Data[34]);
  tran( n15730, Data[35]);
  tran( n15732, Data[36]);
  tran( n15734, Data[37]);
  tran( n15736, Data[38]);
  tran( n15738, Data[39]);
  tran( n15740, Data[40]);
  tran( n15742, Data[41]);
  tran( n15744, Data[42]);
  tran( n15746, Data[43]);
  tran( n15748, Data[44]);
  tran( n15750, Data[45]);
  tran( n15752, Data[46]);
  tran( n15754, Data[47]);
*/
  BUFTD2 \Data_tri[47]  ( .I(n2170), .OE(n2209), .Z(n15754) );
  BUFTD2 \Data_tri[46]  ( .I(n2171), .OE(n2209), .Z(n15752) );
  BUFTD2 \Data_tri[45]  ( .I(n2172), .OE(n2209), .Z(n15750) );
  BUFTD2 \Data_tri[44]  ( .I(n2173), .OE(n2209), .Z(n15748) );
  BUFTD2 \Data_tri[43]  ( .I(n2174), .OE(n2209), .Z(n15746) );
  BUFTD2 \Data_tri[42]  ( .I(n2175), .OE(n2209), .Z(n15744) );
  BUFTD2 \Data_tri[41]  ( .I(n2176), .OE(n2209), .Z(n15742) );
  BUFTD2 \Data_tri[40]  ( .I(n2177), .OE(n2209), .Z(n15740) );
  BUFTD2 \Data_tri[39]  ( .I(n2178), .OE(n2209), .Z(n15738) );
  BUFTD2 \Data_tri[38]  ( .I(n2179), .OE(n2209), .Z(n15736) );
  BUFTD2 \Data_tri[37]  ( .I(n2180), .OE(n2209), .Z(n15734) );
  BUFTD2 \Data_tri[36]  ( .I(n2181), .OE(n2209), .Z(n15732) );
  BUFTD2 \Data_tri[35]  ( .I(n2182), .OE(n2209), .Z(n15730) );
  BUFTD2 \Data_tri[34]  ( .I(n2183), .OE(n2209), .Z(n15728) );
  BUFTD2 \Data_tri[33]  ( .I(n2184), .OE(n2209), .Z(n15726) );
  BUFTD2 \Data_tri[32]  ( .I(n2185), .OE(n2209), .Z(n15724) );
  BUFTD2 \Data_tri[31]  ( .I(n2186), .OE(n2209), .Z(n15722) );
  BUFTD2 \Data_tri[30]  ( .I(n2187), .OE(n2209), .Z(n15720) );
  BUFTD2 \Data_tri[29]  ( .I(n2188), .OE(n2209), .Z(n15718) );
  BUFTD2 \Data_tri[28]  ( .I(n2189), .OE(n2209), .Z(n15716) );
  BUFTD2 \Data_tri[27]  ( .I(n2190), .OE(n2209), .Z(n15714) );
  BUFTD2 \Data_tri[26]  ( .I(n2191), .OE(n2209), .Z(n15712) );
  BUFTD2 \Data_tri[25]  ( .I(n2192), .OE(n2209), .Z(n15710) );
  BUFTD2 \Data_tri[24]  ( .I(n2193), .OE(n2209), .Z(n15708) );
  BUFTD2 \Data_tri[23]  ( .I(n2194), .OE(n2209), .Z(n15706) );
  BUFTD2 \Data_tri[22]  ( .I(n2195), .OE(n2209), .Z(n15704) );
  BUFTD2 \Data_tri[21]  ( .I(n2196), .OE(n2209), .Z(n15702) );
  BUFTD2 \Data_tri[20]  ( .I(n2197), .OE(n2209), .Z(n15700) );
  BUFTD2 \Data_tri[19]  ( .I(n2198), .OE(n2209), .Z(n15698) );
  BUFTD2 \Data_tri[18]  ( .I(n2199), .OE(n2209), .Z(n15696) );
  BUFTD2 \Data_tri[17]  ( .I(n2200), .OE(n2209), .Z(n15694) );
  BUFTD2 \Data_tri[16]  ( .I(n2201), .OE(n2209), .Z(n15692) );
  BUFTD2 \Data_tri[15]  ( .I(n2202), .OE(n2209), .Z(n15690) );
  BUFTD2 \Data_tri[14]  ( .I(n2203), .OE(n2209), .Z(n15688) );
  BUFTD2 \Data_tri[13]  ( .I(n2204), .OE(n2209), .Z(n15686) );
  BUFTD2 \Data_tri[12]  ( .I(n2205), .OE(n2209), .Z(n15684) );
  BUFTD2 \Data_tri[11]  ( .I(n2206), .OE(n2209), .Z(n15682) );
  BUFTD2 \Data_tri[10]  ( .I(n2207), .OE(n2209), .Z(n15680) );
  BUFTD2 \Data_tri[9]  ( .I(n2208), .OE(n2209), .Z(n15678) );
  BUFTD2 \Data_tri[8]  ( .I(n2210), .OE(n2209), .Z(n15676) );
  BUFTD2 \Data_tri[7]  ( .I(n2211), .OE(n2209), .Z(n15674) );
  BUFTD2 \Data_tri[6]  ( .I(n2212), .OE(n2209), .Z(n15672) );
  BUFTD2 \Data_tri[5]  ( .I(n2213), .OE(n2209), .Z(n15670) );
  BUFTD2 \Data_tri[4]  ( .I(n2214), .OE(n2209), .Z(n15668) );
  BUFTD2 \Data_tri[3]  ( .I(n2215), .OE(n2209), .Z(n15666) );
  BUFTD2 \Data_tri[2]  ( .I(n2216), .OE(n2209), .Z(n15664) );
  BUFTD2 \Data_tri[1]  ( .I(n2217), .OE(n2209), .Z(n15662) );
  BUFTD2 \Data_tri[0]  ( .I(n2218), .OE(n2209), .Z(n15660) );
  DFQD1 \Mem_reg[45][47]  ( .D(n6576), .CP(clk), .Q(\Mem[45][47] ) );
  DFQD1 \Mem_reg[45][46]  ( .D(n6574), .CP(clk), .Q(\Mem[45][46] ) );
  DFQD1 \Mem_reg[45][45]  ( .D(n6572), .CP(clk), .Q(\Mem[45][45] ) );
  DFQD1 \Mem_reg[45][44]  ( .D(n6570), .CP(clk), .Q(\Mem[45][44] ) );
  DFQD1 \Mem_reg[45][43]  ( .D(n6568), .CP(clk), .Q(\Mem[45][43] ) );
  DFQD1 \Mem_reg[45][42]  ( .D(n6566), .CP(clk), .Q(\Mem[45][42] ) );
  DFQD1 \Mem_reg[45][41]  ( .D(n6564), .CP(clk), .Q(\Mem[45][41] ) );
  DFQD1 \Mem_reg[45][40]  ( .D(n6562), .CP(clk), .Q(\Mem[45][40] ) );
  DFQD1 \Mem_reg[45][39]  ( .D(n6560), .CP(clk), .Q(\Mem[45][39] ) );
  DFQD1 \Mem_reg[45][38]  ( .D(n6558), .CP(clk), .Q(\Mem[45][38] ) );
  DFQD1 \Mem_reg[45][37]  ( .D(n6556), .CP(clk), .Q(\Mem[45][37] ) );
  DFQD1 \Mem_reg[45][36]  ( .D(n6554), .CP(clk), .Q(\Mem[45][36] ) );
  DFQD1 \Mem_reg[45][35]  ( .D(n6552), .CP(clk), .Q(\Mem[45][35] ) );
  DFQD1 \Mem_reg[45][34]  ( .D(n6550), .CP(clk), .Q(\Mem[45][34] ) );
  DFQD1 \Mem_reg[45][33]  ( .D(n6548), .CP(clk), .Q(\Mem[45][33] ) );
  DFQD1 \Mem_reg[45][32]  ( .D(n6546), .CP(clk), .Q(\Mem[45][32] ) );
  DFQD1 \Mem_reg[45][31]  ( .D(n6544), .CP(clk), .Q(\Mem[45][31] ) );
  DFQD1 \Mem_reg[45][30]  ( .D(n6542), .CP(clk), .Q(\Mem[45][30] ) );
  DFQD1 \Mem_reg[45][29]  ( .D(n6540), .CP(clk), .Q(\Mem[45][29] ) );
  DFQD1 \Mem_reg[45][28]  ( .D(n6538), .CP(clk), .Q(\Mem[45][28] ) );
  DFQD1 \Mem_reg[45][27]  ( .D(n6536), .CP(clk), .Q(\Mem[45][27] ) );
  DFQD1 \Mem_reg[45][26]  ( .D(n6534), .CP(clk), .Q(\Mem[45][26] ) );
  DFQD1 \Mem_reg[45][25]  ( .D(n6532), .CP(clk), .Q(\Mem[45][25] ) );
  DFQD1 \Mem_reg[45][24]  ( .D(n6530), .CP(clk), .Q(\Mem[45][24] ) );
  DFQD1 \Mem_reg[45][23]  ( .D(n6528), .CP(clk), .Q(\Mem[45][23] ) );
  DFQD1 \Mem_reg[45][22]  ( .D(n6526), .CP(clk), .Q(\Mem[45][22] ) );
  DFQD1 \Mem_reg[45][21]  ( .D(n6524), .CP(clk), .Q(\Mem[45][21] ) );
  DFQD1 \Mem_reg[45][20]  ( .D(n6522), .CP(clk), .Q(\Mem[45][20] ) );
  DFQD1 \Mem_reg[45][19]  ( .D(n6520), .CP(clk), .Q(\Mem[45][19] ) );
  DFQD1 \Mem_reg[45][18]  ( .D(n6518), .CP(clk), .Q(\Mem[45][18] ) );
  DFQD1 \Mem_reg[45][17]  ( .D(n6516), .CP(clk), .Q(\Mem[45][17] ) );
  DFQD1 \Mem_reg[45][16]  ( .D(n6514), .CP(clk), .Q(\Mem[45][16] ) );
  DFQD1 \Mem_reg[45][15]  ( .D(n6512), .CP(clk), .Q(\Mem[45][15] ) );
  DFQD1 \Mem_reg[45][14]  ( .D(n6510), .CP(clk), .Q(\Mem[45][14] ) );
  DFQD1 \Mem_reg[45][13]  ( .D(n6508), .CP(clk), .Q(\Mem[45][13] ) );
  DFQD1 \Mem_reg[45][12]  ( .D(n6506), .CP(clk), .Q(\Mem[45][12] ) );
  DFQD1 \Mem_reg[45][11]  ( .D(n6504), .CP(clk), .Q(\Mem[45][11] ) );
  DFQD1 \Mem_reg[45][10]  ( .D(n6502), .CP(clk), .Q(\Mem[45][10] ) );
  DFQD1 \Mem_reg[45][9]  ( .D(n6500), .CP(clk), .Q(\Mem[45][9] ) );
  DFQD1 \Mem_reg[45][8]  ( .D(n6498), .CP(clk), .Q(\Mem[45][8] ) );
  DFQD1 \Mem_reg[45][7]  ( .D(n6496), .CP(clk), .Q(\Mem[45][7] ) );
  DFQD1 \Mem_reg[45][6]  ( .D(n6494), .CP(clk), .Q(\Mem[45][6] ) );
  DFQD1 \Mem_reg[45][5]  ( .D(n6492), .CP(clk), .Q(\Mem[45][5] ) );
  DFQD1 \Mem_reg[45][4]  ( .D(n6490), .CP(clk), .Q(\Mem[45][4] ) );
  DFQD1 \Mem_reg[45][3]  ( .D(n6488), .CP(clk), .Q(\Mem[45][3] ) );
  DFQD1 \Mem_reg[45][2]  ( .D(n6486), .CP(clk), .Q(\Mem[45][2] ) );
  DFQD1 \Mem_reg[45][1]  ( .D(n6484), .CP(clk), .Q(\Mem[45][1] ) );
  DFQD1 \Mem_reg[45][0]  ( .D(n6482), .CP(clk), .Q(\Mem[45][0] ) );
  DFQD1 \Mem_reg[44][47]  ( .D(n6577), .CP(clk), .Q(\Mem[44][47] ) );
  DFQD1 \Mem_reg[44][46]  ( .D(n6575), .CP(clk), .Q(\Mem[44][46] ) );
  DFQD1 \Mem_reg[44][45]  ( .D(n6573), .CP(clk), .Q(\Mem[44][45] ) );
  DFQD1 \Mem_reg[44][44]  ( .D(n6571), .CP(clk), .Q(\Mem[44][44] ) );
  DFQD1 \Mem_reg[44][43]  ( .D(n6569), .CP(clk), .Q(\Mem[44][43] ) );
  DFQD1 \Mem_reg[44][42]  ( .D(n6567), .CP(clk), .Q(\Mem[44][42] ) );
  DFQD1 \Mem_reg[44][41]  ( .D(n6565), .CP(clk), .Q(\Mem[44][41] ) );
  DFQD1 \Mem_reg[44][40]  ( .D(n6563), .CP(clk), .Q(\Mem[44][40] ) );
  DFQD1 \Mem_reg[44][39]  ( .D(n6561), .CP(clk), .Q(\Mem[44][39] ) );
  DFQD1 \Mem_reg[44][38]  ( .D(n6559), .CP(clk), .Q(\Mem[44][38] ) );
  DFQD1 \Mem_reg[44][37]  ( .D(n6557), .CP(clk), .Q(\Mem[44][37] ) );
  DFQD1 \Mem_reg[44][36]  ( .D(n6555), .CP(clk), .Q(\Mem[44][36] ) );
  DFQD1 \Mem_reg[44][35]  ( .D(n6553), .CP(clk), .Q(\Mem[44][35] ) );
  DFQD1 \Mem_reg[44][34]  ( .D(n6551), .CP(clk), .Q(\Mem[44][34] ) );
  DFQD1 \Mem_reg[44][33]  ( .D(n6549), .CP(clk), .Q(\Mem[44][33] ) );
  DFQD1 \Mem_reg[44][32]  ( .D(n6547), .CP(clk), .Q(\Mem[44][32] ) );
  DFQD1 \Mem_reg[44][31]  ( .D(n6545), .CP(clk), .Q(\Mem[44][31] ) );
  DFQD1 \Mem_reg[44][30]  ( .D(n6543), .CP(clk), .Q(\Mem[44][30] ) );
  DFQD1 \Mem_reg[44][29]  ( .D(n6541), .CP(clk), .Q(\Mem[44][29] ) );
  DFQD1 \Mem_reg[44][28]  ( .D(n6539), .CP(clk), .Q(\Mem[44][28] ) );
  DFQD1 \Mem_reg[44][27]  ( .D(n6537), .CP(clk), .Q(\Mem[44][27] ) );
  DFQD1 \Mem_reg[44][26]  ( .D(n6535), .CP(clk), .Q(\Mem[44][26] ) );
  DFQD1 \Mem_reg[44][25]  ( .D(n6533), .CP(clk), .Q(\Mem[44][25] ) );
  DFQD1 \Mem_reg[44][24]  ( .D(n6531), .CP(clk), .Q(\Mem[44][24] ) );
  DFQD1 \Mem_reg[44][23]  ( .D(n6529), .CP(clk), .Q(\Mem[44][23] ) );
  DFQD1 \Mem_reg[44][22]  ( .D(n6527), .CP(clk), .Q(\Mem[44][22] ) );
  DFQD1 \Mem_reg[44][21]  ( .D(n6525), .CP(clk), .Q(\Mem[44][21] ) );
  DFQD1 \Mem_reg[44][20]  ( .D(n6523), .CP(clk), .Q(\Mem[44][20] ) );
  DFQD1 \Mem_reg[44][19]  ( .D(n6521), .CP(clk), .Q(\Mem[44][19] ) );
  DFQD1 \Mem_reg[44][18]  ( .D(n6519), .CP(clk), .Q(\Mem[44][18] ) );
  DFQD1 \Mem_reg[44][17]  ( .D(n6517), .CP(clk), .Q(\Mem[44][17] ) );
  DFQD1 \Mem_reg[44][16]  ( .D(n6515), .CP(clk), .Q(\Mem[44][16] ) );
  DFQD1 \Mem_reg[44][15]  ( .D(n6513), .CP(clk), .Q(\Mem[44][15] ) );
  DFQD1 \Mem_reg[44][14]  ( .D(n6511), .CP(clk), .Q(\Mem[44][14] ) );
  DFQD1 \Mem_reg[44][13]  ( .D(n6509), .CP(clk), .Q(\Mem[44][13] ) );
  DFQD1 \Mem_reg[44][12]  ( .D(n6507), .CP(clk), .Q(\Mem[44][12] ) );
  DFQD1 \Mem_reg[44][11]  ( .D(n6505), .CP(clk), .Q(\Mem[44][11] ) );
  DFQD1 \Mem_reg[44][10]  ( .D(n6503), .CP(clk), .Q(\Mem[44][10] ) );
  DFQD1 \Mem_reg[44][9]  ( .D(n6501), .CP(clk), .Q(\Mem[44][9] ) );
  DFQD1 \Mem_reg[44][8]  ( .D(n6499), .CP(clk), .Q(\Mem[44][8] ) );
  DFQD1 \Mem_reg[44][7]  ( .D(n6497), .CP(clk), .Q(\Mem[44][7] ) );
  DFQD1 \Mem_reg[44][6]  ( .D(n6495), .CP(clk), .Q(\Mem[44][6] ) );
  DFQD1 \Mem_reg[44][5]  ( .D(n6493), .CP(clk), .Q(\Mem[44][5] ) );
  DFQD1 \Mem_reg[44][4]  ( .D(n6491), .CP(clk), .Q(\Mem[44][4] ) );
  DFQD1 \Mem_reg[44][3]  ( .D(n6489), .CP(clk), .Q(\Mem[44][3] ) );
  DFQD1 \Mem_reg[44][2]  ( .D(n6487), .CP(clk), .Q(\Mem[44][2] ) );
  DFQD1 \Mem_reg[44][1]  ( .D(n6485), .CP(clk), .Q(\Mem[44][1] ) );
  DFQD1 \Mem_reg[44][0]  ( .D(n6483), .CP(clk), .Q(\Mem[44][0] ) );
  EDFD1 \Mem_reg[88][47]  ( .D(n24817), .E(n6419), .CP(clk), .Q(n27225) );
  EDFD1 \Mem_reg[87][47]  ( .D(n24817), .E(n6418), .CP(clk), .QN(n6299) );
  EDFD1 \Mem_reg[86][47]  ( .D(n24817), .E(n6417), .CP(clk), .QN(n24700) );
  EDFD1 \Mem_reg[85][47]  ( .D(n24817), .E(n6416), .CP(clk), .QN(n6203) );
  EDFD1 \Mem_reg[84][47]  ( .D(n24817), .E(n6415), .CP(clk), .QN(n6155) );
  EDFD1 \Mem_reg[83][47]  ( .D(n24817), .E(n6414), .CP(clk), .QN(n6107) );
  EDFD1 \Mem_reg[82][47]  ( .D(n24817), .E(n6413), .CP(clk), .QN(n6059) );
  EDFD1 \Mem_reg[81][47]  ( .D(n24817), .E(n6412), .CP(clk), .QN(n6011) );
  EDFD1 \Mem_reg[80][47]  ( .D(n24817), .E(n6411), .CP(clk), .QN(n5963) );
  EDFD1 \Mem_reg[79][47]  ( .D(n24817), .E(n6410), .CP(clk), .QN(n5915) );
  EDFD1 \Mem_reg[78][47]  ( .D(n24817), .E(n6409), .CP(clk), .QN(n5867) );
  EDFD1 \Mem_reg[77][47]  ( .D(n24817), .E(n6408), .CP(clk), .QN(n5819) );
  EDFD1 \Mem_reg[76][47]  ( .D(n24817), .E(n6407), .CP(clk), .QN(n5771) );
  EDFD1 \Mem_reg[75][47]  ( .D(n24817), .E(n6406), .CP(clk), .QN(n27226) );
  EDFD1 \Mem_reg[74][47]  ( .D(n24817), .E(n6405), .CP(clk), .QN(n5675) );
  EDFD1 \Mem_reg[73][47]  ( .D(n24817), .E(n6404), .CP(clk), .QN(n27227) );
  EDFD1 \Mem_reg[72][47]  ( .D(n24817), .E(n6403), .CP(clk), .QN(n5579) );
  EDFD1 \Mem_reg[71][47]  ( .D(n24817), .E(n6402), .CP(clk), .QN(n5531) );
  EDFD1 \Mem_reg[70][47]  ( .D(n24817), .E(n6401), .CP(clk), .QN(n5483) );
  EDFD1 \Mem_reg[69][47]  ( .D(n24817), .E(n6400), .CP(clk), .QN(n5435) );
  EDFD1 \Mem_reg[68][47]  ( .D(n24817), .E(n6399), .CP(clk), .QN(n5387) );
  EDFD1 \Mem_reg[67][47]  ( .D(n24817), .E(n6398), .CP(clk), .QN(n5339) );
  EDFD1 \Mem_reg[66][47]  ( .D(n24817), .E(n6397), .CP(clk), .QN(n5291) );
  EDFD1 \Mem_reg[65][47]  ( .D(n24817), .E(n6396), .CP(clk), .QN(n15637) );
  EDFD1 \Mem_reg[64][47]  ( .D(n24817), .E(n6395), .CP(clk), .QN(n5195) );
  EDFD1 \Mem_reg[63][47]  ( .D(n24817), .E(n6456), .CP(clk), .QN(n5147) );
  EDFD1 \Mem_reg[62][47]  ( .D(n24817), .E(n6455), .CP(clk), .QN(n5099) );
  EDFD1 \Mem_reg[61][47]  ( .D(n24817), .E(n6454), .CP(clk), .QN(n18068) );
  EDFD1 \Mem_reg[60][47]  ( .D(n24817), .E(n6453), .CP(clk), .QN(n18067) );
  EDFD1 \Mem_reg[59][47]  ( .D(n24817), .E(n6452), .CP(clk), .QN(n4955) );
  EDFD1 \Mem_reg[58][47]  ( .D(n24817), .E(n6451), .CP(clk), .QN(n4907) );
  EDFD1 \Mem_reg[57][47]  ( .D(n24817), .E(n6450), .CP(clk), .QN(n4859) );
  EDFD1 \Mem_reg[56][47]  ( .D(n24817), .E(n6449), .CP(clk), .QN(n4811) );
  EDFD1 \Mem_reg[55][47]  ( .D(n24817), .E(n6448), .CP(clk), .QN(n4763) );
  EDFD1 \Mem_reg[54][47]  ( .D(n24817), .E(n6447), .CP(clk), .QN(n15636) );
  EDFD1 \Mem_reg[53][47]  ( .D(n24817), .E(n6446), .CP(clk), .QN(n4667) );
  EDFD1 \Mem_reg[52][47]  ( .D(n24817), .E(n6445), .CP(clk), .Q(n27224) );
  EDFD1 \Mem_reg[51][47]  ( .D(n24817), .E(n6444), .CP(clk), .QN(n4571) );
  EDFD1 \Mem_reg[50][47]  ( .D(n24817), .E(n6443), .CP(clk), .QN(n4523) );
  EDFD1 \Mem_reg[49][47]  ( .D(n24817), .E(n6442), .CP(clk), .QN(n4475) );
  EDFD1 \Mem_reg[48][47]  ( .D(n24817), .E(n6441), .CP(clk), .QN(n4427) );
  EDFD1 \Mem_reg[47][47]  ( .D(n24817), .E(n6440), .CP(clk), .QN(n4379) );
  EDFD1 \Mem_reg[46][47]  ( .D(n24817), .E(n6439), .CP(clk), .QN(n4331) );
  EDFD1 \Mem_reg[43][47]  ( .D(n24817), .E(n6438), .CP(clk), .QN(n4283) );
  EDFD1 \Mem_reg[42][47]  ( .D(n24817), .E(n6437), .CP(clk), .QN(n4235) );
  EDFD1 \Mem_reg[41][47]  ( .D(n24817), .E(n6436), .CP(clk), .QN(n4187) );
  EDFD1 \Mem_reg[40][47]  ( .D(n24817), .E(n6435), .CP(clk), .QN(n4139) );
  EDFD1 \Mem_reg[39][47]  ( .D(n24817), .E(n6434), .CP(clk), .QN(n4091) );
  EDFD1 \Mem_reg[38][47]  ( .D(n24817), .E(n6433), .CP(clk), .QN(n4043) );
  EDFD1 \Mem_reg[37][47]  ( .D(n24817), .E(n6432), .CP(clk), .QN(n3995) );
  EDFD1 \Mem_reg[36][47]  ( .D(n24817), .E(n6431), .CP(clk), .QN(n3947) );
  EDFD1 \Mem_reg[35][47]  ( .D(n24817), .E(n6430), .CP(clk), .QN(n3899) );
  EDFD1 \Mem_reg[34][47]  ( .D(n24817), .E(n6429), .CP(clk), .QN(n3851) );
  EDFD1 \Mem_reg[33][47]  ( .D(n24817), .E(n6428), .CP(clk), .QN(n3803) );
  EDFD1 \Mem_reg[32][47]  ( .D(n24817), .E(n6427), .CP(clk), .QN(n3755) );
  EDFD1 \Mem_reg[31][47]  ( .D(n24817), .E(n6426), .CP(clk), .QN(n3707) );
  EDFD1 \Mem_reg[30][47]  ( .D(n24817), .E(n6425), .CP(clk), .QN(n3659) );
  EDFD1 \Mem_reg[29][47]  ( .D(n24817), .E(n6424), .CP(clk), .QN(n3611) );
  EDFD1 \Mem_reg[28][47]  ( .D(n24817), .E(n6423), .CP(clk), .QN(n3563) );
  EDFD1 \Mem_reg[27][47]  ( .D(n24817), .E(n6422), .CP(clk), .QN(n3515) );
  EDFD1 \Mem_reg[26][47]  ( .D(n24817), .E(n6421), .CP(clk), .QN(n3467) );
  EDFD1 \Mem_reg[25][47]  ( .D(n24817), .E(n6420), .CP(clk), .QN(n3419) );
  EDFD1 \Mem_reg[24][47]  ( .D(n24817), .E(n6463), .CP(clk), .QN(n3371) );
  EDFD1 \Mem_reg[23][47]  ( .D(n24817), .E(n6464), .CP(clk), .QN(n3323) );
  EDFD1 \Mem_reg[22][47]  ( .D(n24817), .E(n6465), .CP(clk), .QN(n3275) );
  EDFD1 \Mem_reg[21][47]  ( .D(n24817), .E(n6466), .CP(clk), .QN(n3227) );
  EDFD1 \Mem_reg[20][47]  ( .D(n24817), .E(n6467), .CP(clk), .QN(n3179) );
  EDFD1 \Mem_reg[19][47]  ( .D(n24817), .E(n6468), .CP(clk), .QN(n3131) );
  EDFD1 \Mem_reg[18][47]  ( .D(n24817), .E(n6469), .CP(clk), .QN(n3083) );
  EDFD1 \Mem_reg[17][47]  ( .D(n24817), .E(n6470), .CP(clk), .QN(n3035) );
  EDFD1 \Mem_reg[16][47]  ( .D(n24817), .E(n6471), .CP(clk), .QN(n2987) );
  EDFD1 \Mem_reg[15][47]  ( .D(n24817), .E(n6472), .CP(clk), .QN(n2939) );
  EDFD1 \Mem_reg[14][47]  ( .D(n24817), .E(n24720), .CP(clk), .QN(n2891) );
  EDFD1 \Mem_reg[13][47]  ( .D(n24817), .E(n24709), .CP(clk), .QN(n2843) );
  EDFD1 \Mem_reg[12][47]  ( .D(n24817), .E(n24717), .CP(clk), .QN(n2795) );
  EDFD1 \Mem_reg[11][47]  ( .D(n24817), .E(n24707), .CP(clk), .QN(n2747) );
  EDFD1 \Mem_reg[10][47]  ( .D(n24817), .E(n6477), .CP(clk), .QN(n2699) );
  EDFD1 \Mem_reg[9][47]  ( .D(n24817), .E(n24708), .CP(clk), .QN(n2651) );
  EDFD1 \Mem_reg[8][47]  ( .D(n24817), .E(n15642), .CP(clk), .QN(n2603) );
  EDFD1 \Mem_reg[7][47]  ( .D(n24817), .E(n24718), .CP(clk), .QN(n2555) );
  EDFD1 \Mem_reg[6][47]  ( .D(n24817), .E(n24716), .CP(clk), .QN(n2507) );
  EDFD1 \Mem_reg[5][47]  ( .D(n24817), .E(n24719), .CP(clk), .QN(n2459) );
  EDFD1 \Mem_reg[4][47]  ( .D(n24817), .E(n24706), .CP(clk), .QN(n2411) );
  EDFD1 \Mem_reg[3][47]  ( .D(n24817), .E(n24721), .CP(clk), .QN(n2363) );
  EDFD1 \Mem_reg[2][47]  ( .D(n24817), .E(n6460), .CP(clk), .QN(n2315) );
  EDFD1 \Mem_reg[1][47]  ( .D(n24817), .E(n24703), .CP(clk), .QN(n2267) );
  EDFD1 \Mem_reg[0][47]  ( .D(n24817), .E(n24705), .CP(clk), .QN(n2219) );
  EDFD1 \Mem_reg[88][46]  ( .D(n24815), .E(n6419), .CP(clk), .Q(n27221) );
  EDFD1 \Mem_reg[87][46]  ( .D(n24815), .E(n6418), .CP(clk), .QN(n6300) );
  EDFD1 \Mem_reg[86][46]  ( .D(n24815), .E(n6417), .CP(clk), .QN(n24697) );
  EDFD1 \Mem_reg[85][46]  ( .D(n24815), .E(n6416), .CP(clk), .QN(n6204) );
  EDFD1 \Mem_reg[84][46]  ( .D(n24815), .E(n6415), .CP(clk), .QN(n6156) );
  EDFD1 \Mem_reg[83][46]  ( .D(n24815), .E(n6414), .CP(clk), .QN(n6108) );
  EDFD1 \Mem_reg[82][46]  ( .D(n24815), .E(n6413), .CP(clk), .QN(n6060) );
  EDFD1 \Mem_reg[81][46]  ( .D(n24815), .E(n6412), .CP(clk), .QN(n6012) );
  EDFD1 \Mem_reg[80][46]  ( .D(n24815), .E(n6411), .CP(clk), .QN(n5964) );
  EDFD1 \Mem_reg[79][46]  ( .D(n24815), .E(n6410), .CP(clk), .QN(n5916) );
  EDFD1 \Mem_reg[78][46]  ( .D(n24815), .E(n6409), .CP(clk), .QN(n5868) );
  EDFD1 \Mem_reg[77][46]  ( .D(n24815), .E(n6408), .CP(clk), .QN(n5820) );
  EDFD1 \Mem_reg[76][46]  ( .D(n24815), .E(n6407), .CP(clk), .QN(n5772) );
  EDFD1 \Mem_reg[75][46]  ( .D(n24815), .E(n6406), .CP(clk), .QN(n27222) );
  EDFD1 \Mem_reg[74][46]  ( .D(n24815), .E(n6405), .CP(clk), .QN(n5676) );
  EDFD1 \Mem_reg[73][46]  ( .D(n24815), .E(n6404), .CP(clk), .QN(n27223) );
  EDFD1 \Mem_reg[72][46]  ( .D(n24815), .E(n6403), .CP(clk), .QN(n5580) );
  EDFD1 \Mem_reg[71][46]  ( .D(n24815), .E(n6402), .CP(clk), .QN(n5532) );
  EDFD1 \Mem_reg[70][46]  ( .D(n24815), .E(n6401), .CP(clk), .QN(n5484) );
  EDFD1 \Mem_reg[69][46]  ( .D(n24815), .E(n6400), .CP(clk), .QN(n5436) );
  EDFD1 \Mem_reg[68][46]  ( .D(n24815), .E(n6399), .CP(clk), .QN(n5388) );
  EDFD1 \Mem_reg[67][46]  ( .D(n24815), .E(n6398), .CP(clk), .QN(n5340) );
  EDFD1 \Mem_reg[66][46]  ( .D(n24815), .E(n6397), .CP(clk), .QN(n5292) );
  EDFD1 \Mem_reg[65][46]  ( .D(n24815), .E(n6396), .CP(clk), .QN(n15633) );
  EDFD1 \Mem_reg[64][46]  ( .D(n24815), .E(n6395), .CP(clk), .QN(n5196) );
  EDFD1 \Mem_reg[63][46]  ( .D(n24815), .E(n6456), .CP(clk), .QN(n5148) );
  EDFD1 \Mem_reg[62][46]  ( .D(n24815), .E(n6455), .CP(clk), .QN(n5100) );
  EDFD1 \Mem_reg[61][46]  ( .D(n24815), .E(n6454), .CP(clk), .QN(n18065) );
  EDFD1 \Mem_reg[60][46]  ( .D(n24815), .E(n6453), .CP(clk), .QN(n18064) );
  EDFD1 \Mem_reg[59][46]  ( .D(n24815), .E(n6452), .CP(clk), .QN(n4956) );
  EDFD1 \Mem_reg[58][46]  ( .D(n24815), .E(n6451), .CP(clk), .QN(n4908) );
  EDFD1 \Mem_reg[57][46]  ( .D(n24815), .E(n6450), .CP(clk), .QN(n4860) );
  EDFD1 \Mem_reg[56][46]  ( .D(n24815), .E(n6449), .CP(clk), .QN(n4812) );
  EDFD1 \Mem_reg[55][46]  ( .D(n24815), .E(n6448), .CP(clk), .QN(n4764) );
  EDFD1 \Mem_reg[54][46]  ( .D(n24815), .E(n6447), .CP(clk), .QN(n15632) );
  EDFD1 \Mem_reg[53][46]  ( .D(n24815), .E(n6446), .CP(clk), .QN(n4668) );
  EDFD1 \Mem_reg[52][46]  ( .D(n24815), .E(n6445), .CP(clk), .Q(n27220) );
  EDFD1 \Mem_reg[51][46]  ( .D(n24815), .E(n6444), .CP(clk), .QN(n4572) );
  EDFD1 \Mem_reg[50][46]  ( .D(n24815), .E(n6443), .CP(clk), .QN(n4524) );
  EDFD1 \Mem_reg[49][46]  ( .D(n24815), .E(n6442), .CP(clk), .QN(n4476) );
  EDFD1 \Mem_reg[48][46]  ( .D(n24815), .E(n6441), .CP(clk), .QN(n4428) );
  EDFD1 \Mem_reg[47][46]  ( .D(n24815), .E(n6440), .CP(clk), .QN(n4380) );
  EDFD1 \Mem_reg[46][46]  ( .D(n24815), .E(n6439), .CP(clk), .QN(n4332) );
  EDFD1 \Mem_reg[43][46]  ( .D(n24815), .E(n6438), .CP(clk), .QN(n4284) );
  EDFD1 \Mem_reg[42][46]  ( .D(n24815), .E(n6437), .CP(clk), .QN(n4236) );
  EDFD1 \Mem_reg[41][46]  ( .D(n24815), .E(n6436), .CP(clk), .QN(n4188) );
  EDFD1 \Mem_reg[40][46]  ( .D(n24815), .E(n6435), .CP(clk), .QN(n4140) );
  EDFD1 \Mem_reg[39][46]  ( .D(n24815), .E(n6434), .CP(clk), .QN(n4092) );
  EDFD1 \Mem_reg[38][46]  ( .D(n24815), .E(n6433), .CP(clk), .QN(n4044) );
  EDFD1 \Mem_reg[37][46]  ( .D(n24815), .E(n6432), .CP(clk), .QN(n3996) );
  EDFD1 \Mem_reg[36][46]  ( .D(n24815), .E(n6431), .CP(clk), .QN(n3948) );
  EDFD1 \Mem_reg[35][46]  ( .D(n24815), .E(n6430), .CP(clk), .QN(n3900) );
  EDFD1 \Mem_reg[34][46]  ( .D(n24815), .E(n6429), .CP(clk), .QN(n3852) );
  EDFD1 \Mem_reg[33][46]  ( .D(n24815), .E(n6428), .CP(clk), .QN(n3804) );
  EDFD1 \Mem_reg[32][46]  ( .D(n24815), .E(n6427), .CP(clk), .QN(n3756) );
  EDFD1 \Mem_reg[31][46]  ( .D(n24815), .E(n6426), .CP(clk), .QN(n3708) );
  EDFD1 \Mem_reg[30][46]  ( .D(n24815), .E(n6425), .CP(clk), .QN(n3660) );
  EDFD1 \Mem_reg[29][46]  ( .D(n24815), .E(n6424), .CP(clk), .QN(n3612) );
  EDFD1 \Mem_reg[28][46]  ( .D(n24815), .E(n6423), .CP(clk), .QN(n3564) );
  EDFD1 \Mem_reg[27][46]  ( .D(n24815), .E(n6422), .CP(clk), .QN(n3516) );
  EDFD1 \Mem_reg[26][46]  ( .D(n24815), .E(n6421), .CP(clk), .QN(n3468) );
  EDFD1 \Mem_reg[25][46]  ( .D(n24815), .E(n6420), .CP(clk), .QN(n3420) );
  EDFD1 \Mem_reg[24][46]  ( .D(n24815), .E(n6463), .CP(clk), .QN(n3372) );
  EDFD1 \Mem_reg[23][46]  ( .D(n24815), .E(n6464), .CP(clk), .QN(n3324) );
  EDFD1 \Mem_reg[22][46]  ( .D(n24815), .E(n6465), .CP(clk), .QN(n3276) );
  EDFD1 \Mem_reg[21][46]  ( .D(n24815), .E(n6466), .CP(clk), .QN(n3228) );
  EDFD1 \Mem_reg[20][46]  ( .D(n24815), .E(n6467), .CP(clk), .QN(n3180) );
  EDFD1 \Mem_reg[19][46]  ( .D(n24815), .E(n6468), .CP(clk), .QN(n3132) );
  EDFD1 \Mem_reg[18][46]  ( .D(n24815), .E(n6469), .CP(clk), .QN(n3084) );
  EDFD1 \Mem_reg[17][46]  ( .D(n24815), .E(n6470), .CP(clk), .QN(n3036) );
  EDFD1 \Mem_reg[16][46]  ( .D(n24815), .E(n6471), .CP(clk), .QN(n2988) );
  EDFD1 \Mem_reg[15][46]  ( .D(n24815), .E(n6472), .CP(clk), .QN(n2940) );
  EDFD1 \Mem_reg[14][46]  ( .D(n24815), .E(n24720), .CP(clk), .QN(n2892) );
  EDFD1 \Mem_reg[13][46]  ( .D(n24815), .E(n24709), .CP(clk), .QN(n2844) );
  EDFD1 \Mem_reg[12][46]  ( .D(n24815), .E(n24717), .CP(clk), .QN(n2796) );
  EDFD1 \Mem_reg[11][46]  ( .D(n24815), .E(n24707), .CP(clk), .QN(n2748) );
  EDFD1 \Mem_reg[10][46]  ( .D(n24815), .E(n6477), .CP(clk), .QN(n2700) );
  EDFD1 \Mem_reg[9][46]  ( .D(n24815), .E(n24708), .CP(clk), .QN(n2652) );
  EDFD1 \Mem_reg[8][46]  ( .D(n24815), .E(n15642), .CP(clk), .QN(n2604) );
  EDFD1 \Mem_reg[7][46]  ( .D(n24815), .E(n24718), .CP(clk), .QN(n2556) );
  EDFD1 \Mem_reg[6][46]  ( .D(n24815), .E(n24716), .CP(clk), .QN(n2508) );
  EDFD1 \Mem_reg[5][46]  ( .D(n24815), .E(n24719), .CP(clk), .QN(n2460) );
  EDFD1 \Mem_reg[4][46]  ( .D(n24815), .E(n24706), .CP(clk), .QN(n2412) );
  EDFD1 \Mem_reg[3][46]  ( .D(n24815), .E(n24721), .CP(clk), .QN(n2364) );
  EDFD1 \Mem_reg[2][46]  ( .D(n24815), .E(n6460), .CP(clk), .QN(n2316) );
  EDFD1 \Mem_reg[1][46]  ( .D(n24815), .E(n24703), .CP(clk), .QN(n2268) );
  EDFD1 \Mem_reg[0][46]  ( .D(n24815), .E(n24705), .CP(clk), .QN(n2220) );
  EDFD1 \Mem_reg[88][45]  ( .D(n24813), .E(n6419), .CP(clk), .Q(n27217) );
  EDFD1 \Mem_reg[87][45]  ( .D(n24813), .E(n6418), .CP(clk), .QN(n6301) );
  EDFD1 \Mem_reg[86][45]  ( .D(n24813), .E(n6417), .CP(clk), .QN(n24694) );
  EDFD1 \Mem_reg[85][45]  ( .D(n24813), .E(n6416), .CP(clk), .QN(n6205) );
  EDFD1 \Mem_reg[84][45]  ( .D(n24813), .E(n6415), .CP(clk), .QN(n6157) );
  EDFD1 \Mem_reg[83][45]  ( .D(n24813), .E(n6414), .CP(clk), .QN(n6109) );
  EDFD1 \Mem_reg[82][45]  ( .D(n24813), .E(n6413), .CP(clk), .QN(n6061) );
  EDFD1 \Mem_reg[81][45]  ( .D(n24813), .E(n6412), .CP(clk), .QN(n6013) );
  EDFD1 \Mem_reg[80][45]  ( .D(n24813), .E(n6411), .CP(clk), .QN(n5965) );
  EDFD1 \Mem_reg[79][45]  ( .D(n24813), .E(n6410), .CP(clk), .QN(n5917) );
  EDFD1 \Mem_reg[78][45]  ( .D(n24813), .E(n6409), .CP(clk), .QN(n5869) );
  EDFD1 \Mem_reg[77][45]  ( .D(n24813), .E(n6408), .CP(clk), .QN(n5821) );
  EDFD1 \Mem_reg[76][45]  ( .D(n24813), .E(n6407), .CP(clk), .QN(n5773) );
  EDFD1 \Mem_reg[75][45]  ( .D(n24813), .E(n6406), .CP(clk), .QN(n27218) );
  EDFD1 \Mem_reg[74][45]  ( .D(n24813), .E(n6405), .CP(clk), .QN(n5677) );
  EDFD1 \Mem_reg[73][45]  ( .D(n24813), .E(n6404), .CP(clk), .QN(n27219) );
  EDFD1 \Mem_reg[72][45]  ( .D(n24813), .E(n6403), .CP(clk), .QN(n5581) );
  EDFD1 \Mem_reg[71][45]  ( .D(n24813), .E(n6402), .CP(clk), .QN(n5533) );
  EDFD1 \Mem_reg[70][45]  ( .D(n24813), .E(n6401), .CP(clk), .QN(n5485) );
  EDFD1 \Mem_reg[69][45]  ( .D(n24813), .E(n6400), .CP(clk), .QN(n5437) );
  EDFD1 \Mem_reg[68][45]  ( .D(n24813), .E(n6399), .CP(clk), .QN(n5389) );
  EDFD1 \Mem_reg[67][45]  ( .D(n24813), .E(n6398), .CP(clk), .QN(n5341) );
  EDFD1 \Mem_reg[66][45]  ( .D(n24813), .E(n6397), .CP(clk), .QN(n5293) );
  EDFD1 \Mem_reg[65][45]  ( .D(n24813), .E(n6396), .CP(clk), .QN(n15629) );
  EDFD1 \Mem_reg[64][45]  ( .D(n24813), .E(n6395), .CP(clk), .QN(n5197) );
  EDFD1 \Mem_reg[63][45]  ( .D(n24813), .E(n6456), .CP(clk), .QN(n5149) );
  EDFD1 \Mem_reg[62][45]  ( .D(n24813), .E(n6455), .CP(clk), .QN(n5101) );
  EDFD1 \Mem_reg[61][45]  ( .D(n24813), .E(n6454), .CP(clk), .QN(n18062) );
  EDFD1 \Mem_reg[60][45]  ( .D(n24813), .E(n6453), .CP(clk), .QN(n18061) );
  EDFD1 \Mem_reg[59][45]  ( .D(n24813), .E(n6452), .CP(clk), .QN(n4957) );
  EDFD1 \Mem_reg[58][45]  ( .D(n24813), .E(n6451), .CP(clk), .QN(n4909) );
  EDFD1 \Mem_reg[57][45]  ( .D(n24813), .E(n6450), .CP(clk), .QN(n4861) );
  EDFD1 \Mem_reg[56][45]  ( .D(n24813), .E(n6449), .CP(clk), .QN(n4813) );
  EDFD1 \Mem_reg[55][45]  ( .D(n24813), .E(n6448), .CP(clk), .QN(n4765) );
  EDFD1 \Mem_reg[54][45]  ( .D(n24813), .E(n6447), .CP(clk), .QN(n15628) );
  EDFD1 \Mem_reg[53][45]  ( .D(n24813), .E(n6446), .CP(clk), .QN(n4669) );
  EDFD1 \Mem_reg[52][45]  ( .D(n24813), .E(n6445), .CP(clk), .Q(n27216) );
  EDFD1 \Mem_reg[51][45]  ( .D(n24813), .E(n6444), .CP(clk), .QN(n4573) );
  EDFD1 \Mem_reg[50][45]  ( .D(n24813), .E(n6443), .CP(clk), .QN(n4525) );
  EDFD1 \Mem_reg[49][45]  ( .D(n24813), .E(n6442), .CP(clk), .QN(n4477) );
  EDFD1 \Mem_reg[48][45]  ( .D(n24813), .E(n6441), .CP(clk), .QN(n4429) );
  EDFD1 \Mem_reg[47][45]  ( .D(n24813), .E(n6440), .CP(clk), .QN(n4381) );
  EDFD1 \Mem_reg[46][45]  ( .D(n24813), .E(n6439), .CP(clk), .QN(n4333) );
  EDFD1 \Mem_reg[43][45]  ( .D(n24813), .E(n6438), .CP(clk), .QN(n4285) );
  EDFD1 \Mem_reg[42][45]  ( .D(n24813), .E(n6437), .CP(clk), .QN(n4237) );
  EDFD1 \Mem_reg[41][45]  ( .D(n24813), .E(n6436), .CP(clk), .QN(n4189) );
  EDFD1 \Mem_reg[40][45]  ( .D(n24813), .E(n6435), .CP(clk), .QN(n4141) );
  EDFD1 \Mem_reg[39][45]  ( .D(n24813), .E(n6434), .CP(clk), .QN(n4093) );
  EDFD1 \Mem_reg[38][45]  ( .D(n24813), .E(n6433), .CP(clk), .QN(n4045) );
  EDFD1 \Mem_reg[37][45]  ( .D(n24813), .E(n6432), .CP(clk), .QN(n3997) );
  EDFD1 \Mem_reg[36][45]  ( .D(n24813), .E(n6431), .CP(clk), .QN(n3949) );
  EDFD1 \Mem_reg[35][45]  ( .D(n24813), .E(n6430), .CP(clk), .QN(n3901) );
  EDFD1 \Mem_reg[34][45]  ( .D(n24813), .E(n6429), .CP(clk), .QN(n3853) );
  EDFD1 \Mem_reg[33][45]  ( .D(n24813), .E(n6428), .CP(clk), .QN(n3805) );
  EDFD1 \Mem_reg[32][45]  ( .D(n24813), .E(n6427), .CP(clk), .QN(n3757) );
  EDFD1 \Mem_reg[31][45]  ( .D(n24813), .E(n6426), .CP(clk), .QN(n3709) );
  EDFD1 \Mem_reg[30][45]  ( .D(n24813), .E(n6425), .CP(clk), .QN(n3661) );
  EDFD1 \Mem_reg[29][45]  ( .D(n24813), .E(n6424), .CP(clk), .QN(n3613) );
  EDFD1 \Mem_reg[28][45]  ( .D(n24813), .E(n6423), .CP(clk), .QN(n3565) );
  EDFD1 \Mem_reg[27][45]  ( .D(n24813), .E(n6422), .CP(clk), .QN(n3517) );
  EDFD1 \Mem_reg[26][45]  ( .D(n24813), .E(n6421), .CP(clk), .QN(n3469) );
  EDFD1 \Mem_reg[25][45]  ( .D(n24813), .E(n6420), .CP(clk), .QN(n3421) );
  EDFD1 \Mem_reg[24][45]  ( .D(n24813), .E(n6463), .CP(clk), .QN(n3373) );
  EDFD1 \Mem_reg[23][45]  ( .D(n24813), .E(n6464), .CP(clk), .QN(n3325) );
  EDFD1 \Mem_reg[22][45]  ( .D(n24813), .E(n6465), .CP(clk), .QN(n3277) );
  EDFD1 \Mem_reg[21][45]  ( .D(n24813), .E(n6466), .CP(clk), .QN(n3229) );
  EDFD1 \Mem_reg[20][45]  ( .D(n24813), .E(n6467), .CP(clk), .QN(n3181) );
  EDFD1 \Mem_reg[19][45]  ( .D(n24813), .E(n6468), .CP(clk), .QN(n3133) );
  EDFD1 \Mem_reg[18][45]  ( .D(n24813), .E(n6469), .CP(clk), .QN(n3085) );
  EDFD1 \Mem_reg[17][45]  ( .D(n24813), .E(n6470), .CP(clk), .QN(n3037) );
  EDFD1 \Mem_reg[16][45]  ( .D(n24813), .E(n6471), .CP(clk), .QN(n2989) );
  EDFD1 \Mem_reg[15][45]  ( .D(n24813), .E(n6472), .CP(clk), .QN(n2941) );
  EDFD1 \Mem_reg[14][45]  ( .D(n24813), .E(n24720), .CP(clk), .QN(n2893) );
  EDFD1 \Mem_reg[13][45]  ( .D(n24813), .E(n24709), .CP(clk), .QN(n2845) );
  EDFD1 \Mem_reg[12][45]  ( .D(n24813), .E(n24717), .CP(clk), .QN(n2797) );
  EDFD1 \Mem_reg[11][45]  ( .D(n24813), .E(n24707), .CP(clk), .QN(n2749) );
  EDFD1 \Mem_reg[10][45]  ( .D(n24813), .E(n6477), .CP(clk), .QN(n2701) );
  EDFD1 \Mem_reg[9][45]  ( .D(n24813), .E(n24708), .CP(clk), .QN(n2653) );
  EDFD1 \Mem_reg[8][45]  ( .D(n24813), .E(n15642), .CP(clk), .QN(n2605) );
  EDFD1 \Mem_reg[7][45]  ( .D(n24813), .E(n24718), .CP(clk), .QN(n2557) );
  EDFD1 \Mem_reg[6][45]  ( .D(n24813), .E(n24716), .CP(clk), .QN(n2509) );
  EDFD1 \Mem_reg[5][45]  ( .D(n24813), .E(n24719), .CP(clk), .QN(n2461) );
  EDFD1 \Mem_reg[4][45]  ( .D(n24813), .E(n24706), .CP(clk), .QN(n2413) );
  EDFD1 \Mem_reg[3][45]  ( .D(n24813), .E(n24721), .CP(clk), .QN(n2365) );
  EDFD1 \Mem_reg[2][45]  ( .D(n24813), .E(n6460), .CP(clk), .QN(n2317) );
  EDFD1 \Mem_reg[1][45]  ( .D(n24813), .E(n24703), .CP(clk), .QN(n2269) );
  EDFD1 \Mem_reg[0][45]  ( .D(n24813), .E(n24705), .CP(clk), .QN(n2221) );
  EDFD1 \Mem_reg[88][44]  ( .D(n24811), .E(n6419), .CP(clk), .Q(n27213) );
  EDFD1 \Mem_reg[87][44]  ( .D(n24811), .E(n6418), .CP(clk), .QN(n6302) );
  EDFD1 \Mem_reg[86][44]  ( .D(n24811), .E(n6417), .CP(clk), .QN(n24691) );
  EDFD1 \Mem_reg[85][44]  ( .D(n24811), .E(n6416), .CP(clk), .QN(n6206) );
  EDFD1 \Mem_reg[84][44]  ( .D(n24811), .E(n6415), .CP(clk), .QN(n6158) );
  EDFD1 \Mem_reg[83][44]  ( .D(n24811), .E(n6414), .CP(clk), .QN(n6110) );
  EDFD1 \Mem_reg[82][44]  ( .D(n24811), .E(n6413), .CP(clk), .QN(n6062) );
  EDFD1 \Mem_reg[81][44]  ( .D(n24811), .E(n6412), .CP(clk), .QN(n6014) );
  EDFD1 \Mem_reg[80][44]  ( .D(n24811), .E(n6411), .CP(clk), .QN(n5966) );
  EDFD1 \Mem_reg[79][44]  ( .D(n24811), .E(n6410), .CP(clk), .QN(n5918) );
  EDFD1 \Mem_reg[78][44]  ( .D(n24811), .E(n6409), .CP(clk), .QN(n5870) );
  EDFD1 \Mem_reg[77][44]  ( .D(n24811), .E(n6408), .CP(clk), .QN(n5822) );
  EDFD1 \Mem_reg[76][44]  ( .D(n24811), .E(n6407), .CP(clk), .QN(n5774) );
  EDFD1 \Mem_reg[75][44]  ( .D(n24811), .E(n6406), .CP(clk), .QN(n27214) );
  EDFD1 \Mem_reg[74][44]  ( .D(n24811), .E(n6405), .CP(clk), .QN(n5678) );
  EDFD1 \Mem_reg[73][44]  ( .D(n24811), .E(n6404), .CP(clk), .QN(n27215) );
  EDFD1 \Mem_reg[72][44]  ( .D(n24811), .E(n6403), .CP(clk), .QN(n5582) );
  EDFD1 \Mem_reg[71][44]  ( .D(n24811), .E(n6402), .CP(clk), .QN(n5534) );
  EDFD1 \Mem_reg[70][44]  ( .D(n24811), .E(n6401), .CP(clk), .QN(n5486) );
  EDFD1 \Mem_reg[69][44]  ( .D(n24811), .E(n6400), .CP(clk), .QN(n5438) );
  EDFD1 \Mem_reg[68][44]  ( .D(n24811), .E(n6399), .CP(clk), .QN(n5390) );
  EDFD1 \Mem_reg[67][44]  ( .D(n24811), .E(n6398), .CP(clk), .QN(n5342) );
  EDFD1 \Mem_reg[66][44]  ( .D(n24811), .E(n6397), .CP(clk), .QN(n5294) );
  EDFD1 \Mem_reg[65][44]  ( .D(n24811), .E(n6396), .CP(clk), .QN(n15625) );
  EDFD1 \Mem_reg[64][44]  ( .D(n24811), .E(n6395), .CP(clk), .QN(n5198) );
  EDFD1 \Mem_reg[63][44]  ( .D(n24811), .E(n6456), .CP(clk), .QN(n5150) );
  EDFD1 \Mem_reg[62][44]  ( .D(n24811), .E(n6455), .CP(clk), .QN(n5102) );
  EDFD1 \Mem_reg[61][44]  ( .D(n24811), .E(n6454), .CP(clk), .QN(n18059) );
  EDFD1 \Mem_reg[60][44]  ( .D(n24811), .E(n6453), .CP(clk), .QN(n18058) );
  EDFD1 \Mem_reg[59][44]  ( .D(n24811), .E(n6452), .CP(clk), .QN(n4958) );
  EDFD1 \Mem_reg[58][44]  ( .D(n24811), .E(n6451), .CP(clk), .QN(n4910) );
  EDFD1 \Mem_reg[57][44]  ( .D(n24811), .E(n6450), .CP(clk), .QN(n4862) );
  EDFD1 \Mem_reg[56][44]  ( .D(n24811), .E(n6449), .CP(clk), .QN(n4814) );
  EDFD1 \Mem_reg[55][44]  ( .D(n24811), .E(n6448), .CP(clk), .QN(n4766) );
  EDFD1 \Mem_reg[54][44]  ( .D(n24811), .E(n6447), .CP(clk), .QN(n15624) );
  EDFD1 \Mem_reg[53][44]  ( .D(n24811), .E(n6446), .CP(clk), .QN(n4670) );
  EDFD1 \Mem_reg[52][44]  ( .D(n24811), .E(n6445), .CP(clk), .Q(n27212) );
  EDFD1 \Mem_reg[51][44]  ( .D(n24811), .E(n6444), .CP(clk), .QN(n4574) );
  EDFD1 \Mem_reg[50][44]  ( .D(n24811), .E(n6443), .CP(clk), .QN(n4526) );
  EDFD1 \Mem_reg[49][44]  ( .D(n24811), .E(n6442), .CP(clk), .QN(n4478) );
  EDFD1 \Mem_reg[48][44]  ( .D(n24811), .E(n6441), .CP(clk), .QN(n4430) );
  EDFD1 \Mem_reg[47][44]  ( .D(n24811), .E(n6440), .CP(clk), .QN(n4382) );
  EDFD1 \Mem_reg[46][44]  ( .D(n24811), .E(n6439), .CP(clk), .QN(n4334) );
  EDFD1 \Mem_reg[43][44]  ( .D(n24811), .E(n6438), .CP(clk), .QN(n4286) );
  EDFD1 \Mem_reg[42][44]  ( .D(n24811), .E(n6437), .CP(clk), .QN(n4238) );
  EDFD1 \Mem_reg[41][44]  ( .D(n24811), .E(n6436), .CP(clk), .QN(n4190) );
  EDFD1 \Mem_reg[40][44]  ( .D(n24811), .E(n6435), .CP(clk), .QN(n4142) );
  EDFD1 \Mem_reg[39][44]  ( .D(n24811), .E(n6434), .CP(clk), .QN(n4094) );
  EDFD1 \Mem_reg[38][44]  ( .D(n24811), .E(n6433), .CP(clk), .QN(n4046) );
  EDFD1 \Mem_reg[37][44]  ( .D(n24811), .E(n6432), .CP(clk), .QN(n3998) );
  EDFD1 \Mem_reg[36][44]  ( .D(n24811), .E(n6431), .CP(clk), .QN(n3950) );
  EDFD1 \Mem_reg[35][44]  ( .D(n24811), .E(n6430), .CP(clk), .QN(n3902) );
  EDFD1 \Mem_reg[34][44]  ( .D(n24811), .E(n6429), .CP(clk), .QN(n3854) );
  EDFD1 \Mem_reg[33][44]  ( .D(n24811), .E(n6428), .CP(clk), .QN(n3806) );
  EDFD1 \Mem_reg[32][44]  ( .D(n24811), .E(n6427), .CP(clk), .QN(n3758) );
  EDFD1 \Mem_reg[31][44]  ( .D(n24811), .E(n6426), .CP(clk), .QN(n3710) );
  EDFD1 \Mem_reg[30][44]  ( .D(n24811), .E(n6425), .CP(clk), .QN(n3662) );
  EDFD1 \Mem_reg[29][44]  ( .D(n24811), .E(n6424), .CP(clk), .QN(n3614) );
  EDFD1 \Mem_reg[28][44]  ( .D(n24811), .E(n6423), .CP(clk), .QN(n3566) );
  EDFD1 \Mem_reg[27][44]  ( .D(n24811), .E(n6422), .CP(clk), .QN(n3518) );
  EDFD1 \Mem_reg[26][44]  ( .D(n24811), .E(n6421), .CP(clk), .QN(n3470) );
  EDFD1 \Mem_reg[25][44]  ( .D(n24811), .E(n6420), .CP(clk), .QN(n3422) );
  EDFD1 \Mem_reg[24][44]  ( .D(n24811), .E(n6463), .CP(clk), .QN(n3374) );
  EDFD1 \Mem_reg[23][44]  ( .D(n24811), .E(n6464), .CP(clk), .QN(n3326) );
  EDFD1 \Mem_reg[22][44]  ( .D(n24811), .E(n6465), .CP(clk), .QN(n3278) );
  EDFD1 \Mem_reg[21][44]  ( .D(n24811), .E(n6466), .CP(clk), .QN(n3230) );
  EDFD1 \Mem_reg[20][44]  ( .D(n24811), .E(n6467), .CP(clk), .QN(n3182) );
  EDFD1 \Mem_reg[19][44]  ( .D(n24811), .E(n6468), .CP(clk), .QN(n3134) );
  EDFD1 \Mem_reg[18][44]  ( .D(n24811), .E(n6469), .CP(clk), .QN(n3086) );
  EDFD1 \Mem_reg[17][44]  ( .D(n24811), .E(n6470), .CP(clk), .QN(n3038) );
  EDFD1 \Mem_reg[16][44]  ( .D(n24811), .E(n6471), .CP(clk), .QN(n2990) );
  EDFD1 \Mem_reg[15][44]  ( .D(n24811), .E(n6472), .CP(clk), .QN(n2942) );
  EDFD1 \Mem_reg[14][44]  ( .D(n24811), .E(n24720), .CP(clk), .QN(n2894) );
  EDFD1 \Mem_reg[13][44]  ( .D(n24811), .E(n24709), .CP(clk), .QN(n2846) );
  EDFD1 \Mem_reg[12][44]  ( .D(n24811), .E(n24717), .CP(clk), .QN(n2798) );
  EDFD1 \Mem_reg[11][44]  ( .D(n24811), .E(n24707), .CP(clk), .QN(n2750) );
  EDFD1 \Mem_reg[10][44]  ( .D(n24811), .E(n6477), .CP(clk), .QN(n2702) );
  EDFD1 \Mem_reg[9][44]  ( .D(n24811), .E(n24708), .CP(clk), .QN(n2654) );
  EDFD1 \Mem_reg[8][44]  ( .D(n24811), .E(n15642), .CP(clk), .QN(n2606) );
  EDFD1 \Mem_reg[7][44]  ( .D(n24811), .E(n24718), .CP(clk), .QN(n2558) );
  EDFD1 \Mem_reg[6][44]  ( .D(n24811), .E(n24716), .CP(clk), .QN(n2510) );
  EDFD1 \Mem_reg[5][44]  ( .D(n24811), .E(n24719), .CP(clk), .QN(n2462) );
  EDFD1 \Mem_reg[4][44]  ( .D(n24811), .E(n24706), .CP(clk), .QN(n2414) );
  EDFD1 \Mem_reg[3][44]  ( .D(n24811), .E(n24721), .CP(clk), .QN(n2366) );
  EDFD1 \Mem_reg[2][44]  ( .D(n24811), .E(n6460), .CP(clk), .QN(n2318) );
  EDFD1 \Mem_reg[1][44]  ( .D(n24811), .E(n24703), .CP(clk), .QN(n2270) );
  EDFD1 \Mem_reg[0][44]  ( .D(n24811), .E(n24705), .CP(clk), .QN(n2222) );
  EDFD1 \Mem_reg[88][43]  ( .D(n24809), .E(n6419), .CP(clk), .Q(n27209) );
  EDFD1 \Mem_reg[87][43]  ( .D(n24809), .E(n6418), .CP(clk), .QN(n6303) );
  EDFD1 \Mem_reg[86][43]  ( .D(n24809), .E(n6417), .CP(clk), .QN(n24688) );
  EDFD1 \Mem_reg[85][43]  ( .D(n24809), .E(n6416), .CP(clk), .QN(n6207) );
  EDFD1 \Mem_reg[84][43]  ( .D(n24809), .E(n6415), .CP(clk), .QN(n6159) );
  EDFD1 \Mem_reg[83][43]  ( .D(n24809), .E(n6414), .CP(clk), .QN(n6111) );
  EDFD1 \Mem_reg[82][43]  ( .D(n24809), .E(n6413), .CP(clk), .QN(n6063) );
  EDFD1 \Mem_reg[81][43]  ( .D(n24809), .E(n6412), .CP(clk), .QN(n6015) );
  EDFD1 \Mem_reg[80][43]  ( .D(n24809), .E(n6411), .CP(clk), .QN(n5967) );
  EDFD1 \Mem_reg[79][43]  ( .D(n24809), .E(n6410), .CP(clk), .QN(n5919) );
  EDFD1 \Mem_reg[78][43]  ( .D(n24809), .E(n6409), .CP(clk), .QN(n5871) );
  EDFD1 \Mem_reg[77][43]  ( .D(n24809), .E(n6408), .CP(clk), .QN(n5823) );
  EDFD1 \Mem_reg[76][43]  ( .D(n24809), .E(n6407), .CP(clk), .QN(n5775) );
  EDFD1 \Mem_reg[75][43]  ( .D(n24809), .E(n6406), .CP(clk), .QN(n27210) );
  EDFD1 \Mem_reg[74][43]  ( .D(n24809), .E(n6405), .CP(clk), .QN(n5679) );
  EDFD1 \Mem_reg[73][43]  ( .D(n24809), .E(n6404), .CP(clk), .QN(n27211) );
  EDFD1 \Mem_reg[72][43]  ( .D(n24809), .E(n6403), .CP(clk), .QN(n5583) );
  EDFD1 \Mem_reg[71][43]  ( .D(n24809), .E(n6402), .CP(clk), .QN(n5535) );
  EDFD1 \Mem_reg[70][43]  ( .D(n24809), .E(n6401), .CP(clk), .QN(n5487) );
  EDFD1 \Mem_reg[69][43]  ( .D(n24809), .E(n6400), .CP(clk), .QN(n5439) );
  EDFD1 \Mem_reg[68][43]  ( .D(n24809), .E(n6399), .CP(clk), .QN(n5391) );
  EDFD1 \Mem_reg[67][43]  ( .D(n24809), .E(n6398), .CP(clk), .QN(n5343) );
  EDFD1 \Mem_reg[66][43]  ( .D(n24809), .E(n6397), .CP(clk), .QN(n5295) );
  EDFD1 \Mem_reg[65][43]  ( .D(n24809), .E(n6396), .CP(clk), .QN(n15621) );
  EDFD1 \Mem_reg[64][43]  ( .D(n24809), .E(n6395), .CP(clk), .QN(n5199) );
  EDFD1 \Mem_reg[63][43]  ( .D(n24809), .E(n6456), .CP(clk), .QN(n5151) );
  EDFD1 \Mem_reg[62][43]  ( .D(n24809), .E(n6455), .CP(clk), .QN(n5103) );
  EDFD1 \Mem_reg[61][43]  ( .D(n24809), .E(n6454), .CP(clk), .QN(n18056) );
  EDFD1 \Mem_reg[60][43]  ( .D(n24809), .E(n6453), .CP(clk), .QN(n18055) );
  EDFD1 \Mem_reg[59][43]  ( .D(n24809), .E(n6452), .CP(clk), .QN(n4959) );
  EDFD1 \Mem_reg[58][43]  ( .D(n24809), .E(n6451), .CP(clk), .QN(n4911) );
  EDFD1 \Mem_reg[57][43]  ( .D(n24809), .E(n6450), .CP(clk), .QN(n4863) );
  EDFD1 \Mem_reg[56][43]  ( .D(n24809), .E(n6449), .CP(clk), .QN(n4815) );
  EDFD1 \Mem_reg[55][43]  ( .D(n24809), .E(n6448), .CP(clk), .QN(n4767) );
  EDFD1 \Mem_reg[54][43]  ( .D(n24809), .E(n6447), .CP(clk), .QN(n15620) );
  EDFD1 \Mem_reg[53][43]  ( .D(n24809), .E(n6446), .CP(clk), .QN(n4671) );
  EDFD1 \Mem_reg[52][43]  ( .D(n24809), .E(n6445), .CP(clk), .Q(n27208) );
  EDFD1 \Mem_reg[51][43]  ( .D(n24809), .E(n6444), .CP(clk), .QN(n4575) );
  EDFD1 \Mem_reg[50][43]  ( .D(n24809), .E(n6443), .CP(clk), .QN(n4527) );
  EDFD1 \Mem_reg[49][43]  ( .D(n24809), .E(n6442), .CP(clk), .QN(n4479) );
  EDFD1 \Mem_reg[48][43]  ( .D(n24809), .E(n6441), .CP(clk), .QN(n4431) );
  EDFD1 \Mem_reg[47][43]  ( .D(n24809), .E(n6440), .CP(clk), .QN(n4383) );
  EDFD1 \Mem_reg[46][43]  ( .D(n24809), .E(n6439), .CP(clk), .QN(n4335) );
  EDFD1 \Mem_reg[43][43]  ( .D(n24809), .E(n6438), .CP(clk), .QN(n4287) );
  EDFD1 \Mem_reg[42][43]  ( .D(n24809), .E(n6437), .CP(clk), .QN(n4239) );
  EDFD1 \Mem_reg[41][43]  ( .D(n24809), .E(n6436), .CP(clk), .QN(n4191) );
  EDFD1 \Mem_reg[40][43]  ( .D(n24809), .E(n6435), .CP(clk), .QN(n4143) );
  EDFD1 \Mem_reg[39][43]  ( .D(n24809), .E(n6434), .CP(clk), .QN(n4095) );
  EDFD1 \Mem_reg[38][43]  ( .D(n24809), .E(n6433), .CP(clk), .QN(n4047) );
  EDFD1 \Mem_reg[37][43]  ( .D(n24809), .E(n6432), .CP(clk), .QN(n3999) );
  EDFD1 \Mem_reg[36][43]  ( .D(n24809), .E(n6431), .CP(clk), .QN(n3951) );
  EDFD1 \Mem_reg[35][43]  ( .D(n24809), .E(n6430), .CP(clk), .QN(n3903) );
  EDFD1 \Mem_reg[34][43]  ( .D(n24809), .E(n6429), .CP(clk), .QN(n3855) );
  EDFD1 \Mem_reg[33][43]  ( .D(n24809), .E(n6428), .CP(clk), .QN(n3807) );
  EDFD1 \Mem_reg[32][43]  ( .D(n24809), .E(n6427), .CP(clk), .QN(n3759) );
  EDFD1 \Mem_reg[31][43]  ( .D(n24809), .E(n6426), .CP(clk), .QN(n3711) );
  EDFD1 \Mem_reg[30][43]  ( .D(n24809), .E(n6425), .CP(clk), .QN(n3663) );
  EDFD1 \Mem_reg[29][43]  ( .D(n24809), .E(n6424), .CP(clk), .QN(n3615) );
  EDFD1 \Mem_reg[28][43]  ( .D(n24809), .E(n6423), .CP(clk), .QN(n3567) );
  EDFD1 \Mem_reg[27][43]  ( .D(n24809), .E(n6422), .CP(clk), .QN(n3519) );
  EDFD1 \Mem_reg[26][43]  ( .D(n24809), .E(n6421), .CP(clk), .QN(n3471) );
  EDFD1 \Mem_reg[25][43]  ( .D(n24809), .E(n6420), .CP(clk), .QN(n3423) );
  EDFD1 \Mem_reg[24][43]  ( .D(n24809), .E(n6463), .CP(clk), .QN(n3375) );
  EDFD1 \Mem_reg[23][43]  ( .D(n24809), .E(n6464), .CP(clk), .QN(n3327) );
  EDFD1 \Mem_reg[22][43]  ( .D(n24809), .E(n6465), .CP(clk), .QN(n3279) );
  EDFD1 \Mem_reg[21][43]  ( .D(n24809), .E(n6466), .CP(clk), .QN(n3231) );
  EDFD1 \Mem_reg[20][43]  ( .D(n24809), .E(n6467), .CP(clk), .QN(n3183) );
  EDFD1 \Mem_reg[19][43]  ( .D(n24809), .E(n6468), .CP(clk), .QN(n3135) );
  EDFD1 \Mem_reg[18][43]  ( .D(n24809), .E(n6469), .CP(clk), .QN(n3087) );
  EDFD1 \Mem_reg[17][43]  ( .D(n24809), .E(n6470), .CP(clk), .QN(n3039) );
  EDFD1 \Mem_reg[16][43]  ( .D(n24809), .E(n6471), .CP(clk), .QN(n2991) );
  EDFD1 \Mem_reg[15][43]  ( .D(n24809), .E(n6472), .CP(clk), .QN(n2943) );
  EDFD1 \Mem_reg[14][43]  ( .D(n24809), .E(n24720), .CP(clk), .QN(n2895) );
  EDFD1 \Mem_reg[13][43]  ( .D(n24809), .E(n24709), .CP(clk), .QN(n2847) );
  EDFD1 \Mem_reg[12][43]  ( .D(n24809), .E(n24717), .CP(clk), .QN(n2799) );
  EDFD1 \Mem_reg[11][43]  ( .D(n24809), .E(n24707), .CP(clk), .QN(n2751) );
  EDFD1 \Mem_reg[10][43]  ( .D(n24809), .E(n6477), .CP(clk), .QN(n2703) );
  EDFD1 \Mem_reg[9][43]  ( .D(n24809), .E(n24708), .CP(clk), .QN(n2655) );
  EDFD1 \Mem_reg[8][43]  ( .D(n24809), .E(n15642), .CP(clk), .QN(n2607) );
  EDFD1 \Mem_reg[7][43]  ( .D(n24809), .E(n24718), .CP(clk), .QN(n2559) );
  EDFD1 \Mem_reg[6][43]  ( .D(n24809), .E(n24716), .CP(clk), .QN(n2511) );
  EDFD1 \Mem_reg[5][43]  ( .D(n24809), .E(n24719), .CP(clk), .QN(n2463) );
  EDFD1 \Mem_reg[4][43]  ( .D(n24809), .E(n24706), .CP(clk), .QN(n2415) );
  EDFD1 \Mem_reg[3][43]  ( .D(n24809), .E(n24721), .CP(clk), .QN(n2367) );
  EDFD1 \Mem_reg[2][43]  ( .D(n24809), .E(n6460), .CP(clk), .QN(n2319) );
  EDFD1 \Mem_reg[1][43]  ( .D(n24809), .E(n24703), .CP(clk), .QN(n2271) );
  EDFD1 \Mem_reg[0][43]  ( .D(n24809), .E(n24705), .CP(clk), .QN(n2223) );
  EDFD1 \Mem_reg[88][42]  ( .D(n24807), .E(n6419), .CP(clk), .Q(n27205) );
  EDFD1 \Mem_reg[87][42]  ( .D(n24807), .E(n6418), .CP(clk), .QN(n6304) );
  EDFD1 \Mem_reg[86][42]  ( .D(n24807), .E(n6417), .CP(clk), .QN(n24685) );
  EDFD1 \Mem_reg[85][42]  ( .D(n24807), .E(n6416), .CP(clk), .QN(n6208) );
  EDFD1 \Mem_reg[84][42]  ( .D(n24807), .E(n6415), .CP(clk), .QN(n6160) );
  EDFD1 \Mem_reg[83][42]  ( .D(n24807), .E(n6414), .CP(clk), .QN(n6112) );
  EDFD1 \Mem_reg[82][42]  ( .D(n24807), .E(n6413), .CP(clk), .QN(n6064) );
  EDFD1 \Mem_reg[81][42]  ( .D(n24807), .E(n6412), .CP(clk), .QN(n6016) );
  EDFD1 \Mem_reg[80][42]  ( .D(n24807), .E(n6411), .CP(clk), .QN(n5968) );
  EDFD1 \Mem_reg[79][42]  ( .D(n24807), .E(n6410), .CP(clk), .QN(n5920) );
  EDFD1 \Mem_reg[78][42]  ( .D(n24807), .E(n6409), .CP(clk), .QN(n5872) );
  EDFD1 \Mem_reg[77][42]  ( .D(n24807), .E(n6408), .CP(clk), .QN(n5824) );
  EDFD1 \Mem_reg[76][42]  ( .D(n24807), .E(n6407), .CP(clk), .QN(n5776) );
  EDFD1 \Mem_reg[75][42]  ( .D(n24807), .E(n6406), .CP(clk), .QN(n27206) );
  EDFD1 \Mem_reg[74][42]  ( .D(n24807), .E(n6405), .CP(clk), .QN(n5680) );
  EDFD1 \Mem_reg[73][42]  ( .D(n24807), .E(n6404), .CP(clk), .QN(n27207) );
  EDFD1 \Mem_reg[72][42]  ( .D(n24807), .E(n6403), .CP(clk), .QN(n5584) );
  EDFD1 \Mem_reg[71][42]  ( .D(n24807), .E(n6402), .CP(clk), .QN(n5536) );
  EDFD1 \Mem_reg[70][42]  ( .D(n24807), .E(n6401), .CP(clk), .QN(n5488) );
  EDFD1 \Mem_reg[69][42]  ( .D(n24807), .E(n6400), .CP(clk), .QN(n5440) );
  EDFD1 \Mem_reg[68][42]  ( .D(n24807), .E(n6399), .CP(clk), .QN(n5392) );
  EDFD1 \Mem_reg[67][42]  ( .D(n24807), .E(n6398), .CP(clk), .QN(n5344) );
  EDFD1 \Mem_reg[66][42]  ( .D(n24807), .E(n6397), .CP(clk), .QN(n5296) );
  EDFD1 \Mem_reg[65][42]  ( .D(n24807), .E(n6396), .CP(clk), .QN(n15617) );
  EDFD1 \Mem_reg[64][42]  ( .D(n24807), .E(n6395), .CP(clk), .QN(n5200) );
  EDFD1 \Mem_reg[63][42]  ( .D(n24807), .E(n6456), .CP(clk), .QN(n5152) );
  EDFD1 \Mem_reg[62][42]  ( .D(n24807), .E(n6455), .CP(clk), .QN(n5104) );
  EDFD1 \Mem_reg[61][42]  ( .D(n24807), .E(n6454), .CP(clk), .QN(n18053) );
  EDFD1 \Mem_reg[60][42]  ( .D(n24807), .E(n6453), .CP(clk), .QN(n18052) );
  EDFD1 \Mem_reg[59][42]  ( .D(n24807), .E(n6452), .CP(clk), .QN(n4960) );
  EDFD1 \Mem_reg[58][42]  ( .D(n24807), .E(n6451), .CP(clk), .QN(n4912) );
  EDFD1 \Mem_reg[57][42]  ( .D(n24807), .E(n6450), .CP(clk), .QN(n4864) );
  EDFD1 \Mem_reg[56][42]  ( .D(n24807), .E(n6449), .CP(clk), .QN(n4816) );
  EDFD1 \Mem_reg[55][42]  ( .D(n24807), .E(n6448), .CP(clk), .QN(n4768) );
  EDFD1 \Mem_reg[54][42]  ( .D(n24807), .E(n6447), .CP(clk), .QN(n15616) );
  EDFD1 \Mem_reg[53][42]  ( .D(n24807), .E(n6446), .CP(clk), .QN(n4672) );
  EDFD1 \Mem_reg[52][42]  ( .D(n24807), .E(n6445), .CP(clk), .Q(n27204) );
  EDFD1 \Mem_reg[51][42]  ( .D(n24807), .E(n6444), .CP(clk), .QN(n4576) );
  EDFD1 \Mem_reg[50][42]  ( .D(n24807), .E(n6443), .CP(clk), .QN(n4528) );
  EDFD1 \Mem_reg[49][42]  ( .D(n24807), .E(n6442), .CP(clk), .QN(n4480) );
  EDFD1 \Mem_reg[48][42]  ( .D(n24807), .E(n6441), .CP(clk), .QN(n4432) );
  EDFD1 \Mem_reg[47][42]  ( .D(n24807), .E(n6440), .CP(clk), .QN(n4384) );
  EDFD1 \Mem_reg[46][42]  ( .D(n24807), .E(n6439), .CP(clk), .QN(n4336) );
  EDFD1 \Mem_reg[43][42]  ( .D(n24807), .E(n6438), .CP(clk), .QN(n4288) );
  EDFD1 \Mem_reg[42][42]  ( .D(n24807), .E(n6437), .CP(clk), .QN(n4240) );
  EDFD1 \Mem_reg[41][42]  ( .D(n24807), .E(n6436), .CP(clk), .QN(n4192) );
  EDFD1 \Mem_reg[40][42]  ( .D(n24807), .E(n6435), .CP(clk), .QN(n4144) );
  EDFD1 \Mem_reg[39][42]  ( .D(n24807), .E(n6434), .CP(clk), .QN(n4096) );
  EDFD1 \Mem_reg[38][42]  ( .D(n24807), .E(n6433), .CP(clk), .QN(n4048) );
  EDFD1 \Mem_reg[37][42]  ( .D(n24807), .E(n6432), .CP(clk), .QN(n4000) );
  EDFD1 \Mem_reg[36][42]  ( .D(n24807), .E(n6431), .CP(clk), .QN(n3952) );
  EDFD1 \Mem_reg[35][42]  ( .D(n24807), .E(n6430), .CP(clk), .QN(n3904) );
  EDFD1 \Mem_reg[34][42]  ( .D(n24807), .E(n6429), .CP(clk), .QN(n3856) );
  EDFD1 \Mem_reg[33][42]  ( .D(n24807), .E(n6428), .CP(clk), .QN(n3808) );
  EDFD1 \Mem_reg[32][42]  ( .D(n24807), .E(n6427), .CP(clk), .QN(n3760) );
  EDFD1 \Mem_reg[31][42]  ( .D(n24807), .E(n6426), .CP(clk), .QN(n3712) );
  EDFD1 \Mem_reg[30][42]  ( .D(n24807), .E(n6425), .CP(clk), .QN(n3664) );
  EDFD1 \Mem_reg[29][42]  ( .D(n24807), .E(n6424), .CP(clk), .QN(n3616) );
  EDFD1 \Mem_reg[28][42]  ( .D(n24807), .E(n6423), .CP(clk), .QN(n3568) );
  EDFD1 \Mem_reg[27][42]  ( .D(n24807), .E(n6422), .CP(clk), .QN(n3520) );
  EDFD1 \Mem_reg[26][42]  ( .D(n24807), .E(n6421), .CP(clk), .QN(n3472) );
  EDFD1 \Mem_reg[25][42]  ( .D(n24807), .E(n6420), .CP(clk), .QN(n3424) );
  EDFD1 \Mem_reg[24][42]  ( .D(n24807), .E(n6463), .CP(clk), .QN(n3376) );
  EDFD1 \Mem_reg[23][42]  ( .D(n24807), .E(n6464), .CP(clk), .QN(n3328) );
  EDFD1 \Mem_reg[22][42]  ( .D(n24807), .E(n6465), .CP(clk), .QN(n3280) );
  EDFD1 \Mem_reg[21][42]  ( .D(n24807), .E(n6466), .CP(clk), .QN(n3232) );
  EDFD1 \Mem_reg[20][42]  ( .D(n24807), .E(n6467), .CP(clk), .QN(n3184) );
  EDFD1 \Mem_reg[19][42]  ( .D(n24807), .E(n6468), .CP(clk), .QN(n3136) );
  EDFD1 \Mem_reg[18][42]  ( .D(n24807), .E(n6469), .CP(clk), .QN(n3088) );
  EDFD1 \Mem_reg[17][42]  ( .D(n24807), .E(n6470), .CP(clk), .QN(n3040) );
  EDFD1 \Mem_reg[16][42]  ( .D(n24807), .E(n6471), .CP(clk), .QN(n2992) );
  EDFD1 \Mem_reg[15][42]  ( .D(n24807), .E(n6472), .CP(clk), .QN(n2944) );
  EDFD1 \Mem_reg[14][42]  ( .D(n24807), .E(n24720), .CP(clk), .QN(n2896) );
  EDFD1 \Mem_reg[13][42]  ( .D(n24807), .E(n24709), .CP(clk), .QN(n2848) );
  EDFD1 \Mem_reg[12][42]  ( .D(n24807), .E(n24717), .CP(clk), .QN(n2800) );
  EDFD1 \Mem_reg[11][42]  ( .D(n24807), .E(n24707), .CP(clk), .QN(n2752) );
  EDFD1 \Mem_reg[10][42]  ( .D(n24807), .E(n6477), .CP(clk), .QN(n2704) );
  EDFD1 \Mem_reg[9][42]  ( .D(n24807), .E(n24708), .CP(clk), .QN(n2656) );
  EDFD1 \Mem_reg[8][42]  ( .D(n24807), .E(n15642), .CP(clk), .QN(n2608) );
  EDFD1 \Mem_reg[7][42]  ( .D(n24807), .E(n24718), .CP(clk), .QN(n2560) );
  EDFD1 \Mem_reg[6][42]  ( .D(n24807), .E(n24716), .CP(clk), .QN(n2512) );
  EDFD1 \Mem_reg[5][42]  ( .D(n24807), .E(n24719), .CP(clk), .QN(n2464) );
  EDFD1 \Mem_reg[4][42]  ( .D(n24807), .E(n24706), .CP(clk), .QN(n2416) );
  EDFD1 \Mem_reg[3][42]  ( .D(n24807), .E(n24721), .CP(clk), .QN(n2368) );
  EDFD1 \Mem_reg[2][42]  ( .D(n24807), .E(n6460), .CP(clk), .QN(n2320) );
  EDFD1 \Mem_reg[1][42]  ( .D(n24807), .E(n24703), .CP(clk), .QN(n2272) );
  EDFD1 \Mem_reg[0][42]  ( .D(n24807), .E(n24705), .CP(clk), .QN(n2224) );
  EDFD1 \Mem_reg[88][41]  ( .D(n24805), .E(n6419), .CP(clk), .Q(n27201) );
  EDFD1 \Mem_reg[87][41]  ( .D(n24805), .E(n6418), .CP(clk), .QN(n6305) );
  EDFD1 \Mem_reg[86][41]  ( .D(n24805), .E(n6417), .CP(clk), .QN(n24682) );
  EDFD1 \Mem_reg[85][41]  ( .D(n24805), .E(n6416), .CP(clk), .QN(n6209) );
  EDFD1 \Mem_reg[84][41]  ( .D(n24805), .E(n6415), .CP(clk), .QN(n6161) );
  EDFD1 \Mem_reg[83][41]  ( .D(n24805), .E(n6414), .CP(clk), .QN(n6113) );
  EDFD1 \Mem_reg[82][41]  ( .D(n24805), .E(n6413), .CP(clk), .QN(n6065) );
  EDFD1 \Mem_reg[81][41]  ( .D(n24805), .E(n6412), .CP(clk), .QN(n6017) );
  EDFD1 \Mem_reg[80][41]  ( .D(n24805), .E(n6411), .CP(clk), .QN(n5969) );
  EDFD1 \Mem_reg[79][41]  ( .D(n24805), .E(n6410), .CP(clk), .QN(n5921) );
  EDFD1 \Mem_reg[78][41]  ( .D(n24805), .E(n6409), .CP(clk), .QN(n5873) );
  EDFD1 \Mem_reg[77][41]  ( .D(n24805), .E(n6408), .CP(clk), .QN(n5825) );
  EDFD1 \Mem_reg[76][41]  ( .D(n24805), .E(n6407), .CP(clk), .QN(n5777) );
  EDFD1 \Mem_reg[75][41]  ( .D(n24805), .E(n6406), .CP(clk), .QN(n27202) );
  EDFD1 \Mem_reg[74][41]  ( .D(n24805), .E(n6405), .CP(clk), .QN(n5681) );
  EDFD1 \Mem_reg[73][41]  ( .D(n24805), .E(n6404), .CP(clk), .QN(n27203) );
  EDFD1 \Mem_reg[72][41]  ( .D(n24805), .E(n6403), .CP(clk), .QN(n5585) );
  EDFD1 \Mem_reg[71][41]  ( .D(n24805), .E(n6402), .CP(clk), .QN(n5537) );
  EDFD1 \Mem_reg[70][41]  ( .D(n24805), .E(n6401), .CP(clk), .QN(n5489) );
  EDFD1 \Mem_reg[69][41]  ( .D(n24805), .E(n6400), .CP(clk), .QN(n5441) );
  EDFD1 \Mem_reg[68][41]  ( .D(n24805), .E(n6399), .CP(clk), .QN(n5393) );
  EDFD1 \Mem_reg[67][41]  ( .D(n24805), .E(n6398), .CP(clk), .QN(n5345) );
  EDFD1 \Mem_reg[66][41]  ( .D(n24805), .E(n6397), .CP(clk), .QN(n5297) );
  EDFD1 \Mem_reg[65][41]  ( .D(n24805), .E(n6396), .CP(clk), .QN(n15613) );
  EDFD1 \Mem_reg[64][41]  ( .D(n24805), .E(n6395), .CP(clk), .QN(n5201) );
  EDFD1 \Mem_reg[63][41]  ( .D(n24805), .E(n6456), .CP(clk), .QN(n5153) );
  EDFD1 \Mem_reg[62][41]  ( .D(n24805), .E(n6455), .CP(clk), .QN(n5105) );
  EDFD1 \Mem_reg[61][41]  ( .D(n24805), .E(n6454), .CP(clk), .QN(n18050) );
  EDFD1 \Mem_reg[60][41]  ( .D(n24805), .E(n6453), .CP(clk), .QN(n18049) );
  EDFD1 \Mem_reg[59][41]  ( .D(n24805), .E(n6452), .CP(clk), .QN(n4961) );
  EDFD1 \Mem_reg[58][41]  ( .D(n24805), .E(n6451), .CP(clk), .QN(n4913) );
  EDFD1 \Mem_reg[57][41]  ( .D(n24805), .E(n6450), .CP(clk), .QN(n4865) );
  EDFD1 \Mem_reg[56][41]  ( .D(n24805), .E(n6449), .CP(clk), .QN(n4817) );
  EDFD1 \Mem_reg[55][41]  ( .D(n24805), .E(n6448), .CP(clk), .QN(n4769) );
  EDFD1 \Mem_reg[54][41]  ( .D(n24805), .E(n6447), .CP(clk), .QN(n15612) );
  EDFD1 \Mem_reg[53][41]  ( .D(n24805), .E(n6446), .CP(clk), .QN(n4673) );
  EDFD1 \Mem_reg[52][41]  ( .D(n24805), .E(n6445), .CP(clk), .Q(n27200) );
  EDFD1 \Mem_reg[51][41]  ( .D(n24805), .E(n6444), .CP(clk), .QN(n4577) );
  EDFD1 \Mem_reg[50][41]  ( .D(n24805), .E(n6443), .CP(clk), .QN(n4529) );
  EDFD1 \Mem_reg[49][41]  ( .D(n24805), .E(n6442), .CP(clk), .QN(n4481) );
  EDFD1 \Mem_reg[48][41]  ( .D(n24805), .E(n6441), .CP(clk), .QN(n4433) );
  EDFD1 \Mem_reg[47][41]  ( .D(n24805), .E(n6440), .CP(clk), .QN(n4385) );
  EDFD1 \Mem_reg[46][41]  ( .D(n24805), .E(n6439), .CP(clk), .QN(n4337) );
  EDFD1 \Mem_reg[43][41]  ( .D(n24805), .E(n6438), .CP(clk), .QN(n4289) );
  EDFD1 \Mem_reg[42][41]  ( .D(n24805), .E(n6437), .CP(clk), .QN(n4241) );
  EDFD1 \Mem_reg[41][41]  ( .D(n24805), .E(n6436), .CP(clk), .QN(n4193) );
  EDFD1 \Mem_reg[40][41]  ( .D(n24805), .E(n6435), .CP(clk), .QN(n4145) );
  EDFD1 \Mem_reg[39][41]  ( .D(n24805), .E(n6434), .CP(clk), .QN(n4097) );
  EDFD1 \Mem_reg[38][41]  ( .D(n24805), .E(n6433), .CP(clk), .QN(n4049) );
  EDFD1 \Mem_reg[37][41]  ( .D(n24805), .E(n6432), .CP(clk), .QN(n4001) );
  EDFD1 \Mem_reg[36][41]  ( .D(n24805), .E(n6431), .CP(clk), .QN(n3953) );
  EDFD1 \Mem_reg[35][41]  ( .D(n24805), .E(n6430), .CP(clk), .QN(n3905) );
  EDFD1 \Mem_reg[34][41]  ( .D(n24805), .E(n6429), .CP(clk), .QN(n3857) );
  EDFD1 \Mem_reg[33][41]  ( .D(n24805), .E(n6428), .CP(clk), .QN(n3809) );
  EDFD1 \Mem_reg[32][41]  ( .D(n24805), .E(n6427), .CP(clk), .QN(n3761) );
  EDFD1 \Mem_reg[31][41]  ( .D(n24805), .E(n6426), .CP(clk), .QN(n3713) );
  EDFD1 \Mem_reg[30][41]  ( .D(n24805), .E(n6425), .CP(clk), .QN(n3665) );
  EDFD1 \Mem_reg[29][41]  ( .D(n24805), .E(n6424), .CP(clk), .QN(n3617) );
  EDFD1 \Mem_reg[28][41]  ( .D(n24805), .E(n6423), .CP(clk), .QN(n3569) );
  EDFD1 \Mem_reg[27][41]  ( .D(n24805), .E(n6422), .CP(clk), .QN(n3521) );
  EDFD1 \Mem_reg[26][41]  ( .D(n24805), .E(n6421), .CP(clk), .QN(n3473) );
  EDFD1 \Mem_reg[25][41]  ( .D(n24805), .E(n6420), .CP(clk), .QN(n3425) );
  EDFD1 \Mem_reg[24][41]  ( .D(n24805), .E(n6463), .CP(clk), .QN(n3377) );
  EDFD1 \Mem_reg[23][41]  ( .D(n24805), .E(n6464), .CP(clk), .QN(n3329) );
  EDFD1 \Mem_reg[22][41]  ( .D(n24805), .E(n6465), .CP(clk), .QN(n3281) );
  EDFD1 \Mem_reg[21][41]  ( .D(n24805), .E(n6466), .CP(clk), .QN(n3233) );
  EDFD1 \Mem_reg[20][41]  ( .D(n24805), .E(n6467), .CP(clk), .QN(n3185) );
  EDFD1 \Mem_reg[19][41]  ( .D(n24805), .E(n6468), .CP(clk), .QN(n3137) );
  EDFD1 \Mem_reg[18][41]  ( .D(n24805), .E(n6469), .CP(clk), .QN(n3089) );
  EDFD1 \Mem_reg[17][41]  ( .D(n24805), .E(n6470), .CP(clk), .QN(n3041) );
  EDFD1 \Mem_reg[16][41]  ( .D(n24805), .E(n6471), .CP(clk), .QN(n2993) );
  EDFD1 \Mem_reg[15][41]  ( .D(n24805), .E(n6472), .CP(clk), .QN(n2945) );
  EDFD1 \Mem_reg[14][41]  ( .D(n24805), .E(n24720), .CP(clk), .QN(n2897) );
  EDFD1 \Mem_reg[13][41]  ( .D(n24805), .E(n24709), .CP(clk), .QN(n2849) );
  EDFD1 \Mem_reg[12][41]  ( .D(n24805), .E(n24717), .CP(clk), .QN(n2801) );
  EDFD1 \Mem_reg[11][41]  ( .D(n24805), .E(n24707), .CP(clk), .QN(n2753) );
  EDFD1 \Mem_reg[10][41]  ( .D(n24805), .E(n6477), .CP(clk), .QN(n2705) );
  EDFD1 \Mem_reg[9][41]  ( .D(n24805), .E(n24708), .CP(clk), .QN(n2657) );
  EDFD1 \Mem_reg[8][41]  ( .D(n24805), .E(n15642), .CP(clk), .QN(n2609) );
  EDFD1 \Mem_reg[7][41]  ( .D(n24805), .E(n24718), .CP(clk), .QN(n2561) );
  EDFD1 \Mem_reg[6][41]  ( .D(n24805), .E(n24716), .CP(clk), .QN(n2513) );
  EDFD1 \Mem_reg[5][41]  ( .D(n24805), .E(n24719), .CP(clk), .QN(n2465) );
  EDFD1 \Mem_reg[4][41]  ( .D(n24805), .E(n24706), .CP(clk), .QN(n2417) );
  EDFD1 \Mem_reg[3][41]  ( .D(n24805), .E(n24721), .CP(clk), .QN(n2369) );
  EDFD1 \Mem_reg[2][41]  ( .D(n24805), .E(n6460), .CP(clk), .QN(n2321) );
  EDFD1 \Mem_reg[1][41]  ( .D(n24805), .E(n24703), .CP(clk), .QN(n2273) );
  EDFD1 \Mem_reg[0][41]  ( .D(n24805), .E(n24705), .CP(clk), .QN(n2225) );
  EDFD1 \Mem_reg[88][40]  ( .D(n24803), .E(n6419), .CP(clk), .Q(n27197) );
  EDFD1 \Mem_reg[87][40]  ( .D(n24803), .E(n6418), .CP(clk), .QN(n6306) );
  EDFD1 \Mem_reg[86][40]  ( .D(n24803), .E(n6417), .CP(clk), .QN(n24679) );
  EDFD1 \Mem_reg[85][40]  ( .D(n24803), .E(n6416), .CP(clk), .QN(n6210) );
  EDFD1 \Mem_reg[84][40]  ( .D(n24803), .E(n6415), .CP(clk), .QN(n6162) );
  EDFD1 \Mem_reg[83][40]  ( .D(n24803), .E(n6414), .CP(clk), .QN(n6114) );
  EDFD1 \Mem_reg[82][40]  ( .D(n24803), .E(n6413), .CP(clk), .QN(n6066) );
  EDFD1 \Mem_reg[81][40]  ( .D(n24803), .E(n6412), .CP(clk), .QN(n6018) );
  EDFD1 \Mem_reg[80][40]  ( .D(n24803), .E(n6411), .CP(clk), .QN(n5970) );
  EDFD1 \Mem_reg[79][40]  ( .D(n24803), .E(n6410), .CP(clk), .QN(n5922) );
  EDFD1 \Mem_reg[78][40]  ( .D(n24803), .E(n6409), .CP(clk), .QN(n5874) );
  EDFD1 \Mem_reg[77][40]  ( .D(n24803), .E(n6408), .CP(clk), .QN(n5826) );
  EDFD1 \Mem_reg[76][40]  ( .D(n24803), .E(n6407), .CP(clk), .QN(n5778) );
  EDFD1 \Mem_reg[75][40]  ( .D(n24803), .E(n6406), .CP(clk), .QN(n27198) );
  EDFD1 \Mem_reg[74][40]  ( .D(n24803), .E(n6405), .CP(clk), .QN(n5682) );
  EDFD1 \Mem_reg[73][40]  ( .D(n24803), .E(n6404), .CP(clk), .QN(n27199) );
  EDFD1 \Mem_reg[72][40]  ( .D(n24803), .E(n6403), .CP(clk), .QN(n5586) );
  EDFD1 \Mem_reg[71][40]  ( .D(n24803), .E(n6402), .CP(clk), .QN(n5538) );
  EDFD1 \Mem_reg[70][40]  ( .D(n24803), .E(n6401), .CP(clk), .QN(n5490) );
  EDFD1 \Mem_reg[69][40]  ( .D(n24803), .E(n6400), .CP(clk), .QN(n5442) );
  EDFD1 \Mem_reg[68][40]  ( .D(n24803), .E(n6399), .CP(clk), .QN(n5394) );
  EDFD1 \Mem_reg[67][40]  ( .D(n24803), .E(n6398), .CP(clk), .QN(n5346) );
  EDFD1 \Mem_reg[66][40]  ( .D(n24803), .E(n6397), .CP(clk), .QN(n5298) );
  EDFD1 \Mem_reg[65][40]  ( .D(n24803), .E(n6396), .CP(clk), .QN(n15609) );
  EDFD1 \Mem_reg[64][40]  ( .D(n24803), .E(n6395), .CP(clk), .QN(n5202) );
  EDFD1 \Mem_reg[63][40]  ( .D(n24803), .E(n6456), .CP(clk), .QN(n5154) );
  EDFD1 \Mem_reg[62][40]  ( .D(n24803), .E(n6455), .CP(clk), .QN(n5106) );
  EDFD1 \Mem_reg[61][40]  ( .D(n24803), .E(n6454), .CP(clk), .QN(n18047) );
  EDFD1 \Mem_reg[60][40]  ( .D(n24803), .E(n6453), .CP(clk), .QN(n18046) );
  EDFD1 \Mem_reg[59][40]  ( .D(n24803), .E(n6452), .CP(clk), .QN(n4962) );
  EDFD1 \Mem_reg[58][40]  ( .D(n24803), .E(n6451), .CP(clk), .QN(n4914) );
  EDFD1 \Mem_reg[57][40]  ( .D(n24803), .E(n6450), .CP(clk), .QN(n4866) );
  EDFD1 \Mem_reg[56][40]  ( .D(n24803), .E(n6449), .CP(clk), .QN(n4818) );
  EDFD1 \Mem_reg[55][40]  ( .D(n24803), .E(n6448), .CP(clk), .QN(n4770) );
  EDFD1 \Mem_reg[54][40]  ( .D(n24803), .E(n6447), .CP(clk), .QN(n15608) );
  EDFD1 \Mem_reg[53][40]  ( .D(n24803), .E(n6446), .CP(clk), .QN(n4674) );
  EDFD1 \Mem_reg[52][40]  ( .D(n24803), .E(n6445), .CP(clk), .Q(n27196) );
  EDFD1 \Mem_reg[51][40]  ( .D(n24803), .E(n6444), .CP(clk), .QN(n4578) );
  EDFD1 \Mem_reg[50][40]  ( .D(n24803), .E(n6443), .CP(clk), .QN(n4530) );
  EDFD1 \Mem_reg[49][40]  ( .D(n24803), .E(n6442), .CP(clk), .QN(n4482) );
  EDFD1 \Mem_reg[48][40]  ( .D(n24803), .E(n6441), .CP(clk), .QN(n4434) );
  EDFD1 \Mem_reg[47][40]  ( .D(n24803), .E(n6440), .CP(clk), .QN(n4386) );
  EDFD1 \Mem_reg[46][40]  ( .D(n24803), .E(n6439), .CP(clk), .QN(n4338) );
  EDFD1 \Mem_reg[43][40]  ( .D(n24803), .E(n6438), .CP(clk), .QN(n4290) );
  EDFD1 \Mem_reg[42][40]  ( .D(n24803), .E(n6437), .CP(clk), .QN(n4242) );
  EDFD1 \Mem_reg[41][40]  ( .D(n24803), .E(n6436), .CP(clk), .QN(n4194) );
  EDFD1 \Mem_reg[40][40]  ( .D(n24803), .E(n6435), .CP(clk), .QN(n4146) );
  EDFD1 \Mem_reg[39][40]  ( .D(n24803), .E(n6434), .CP(clk), .QN(n4098) );
  EDFD1 \Mem_reg[38][40]  ( .D(n24803), .E(n6433), .CP(clk), .QN(n4050) );
  EDFD1 \Mem_reg[37][40]  ( .D(n24803), .E(n6432), .CP(clk), .QN(n4002) );
  EDFD1 \Mem_reg[36][40]  ( .D(n24803), .E(n6431), .CP(clk), .QN(n3954) );
  EDFD1 \Mem_reg[35][40]  ( .D(n24803), .E(n6430), .CP(clk), .QN(n3906) );
  EDFD1 \Mem_reg[34][40]  ( .D(n24803), .E(n6429), .CP(clk), .QN(n3858) );
  EDFD1 \Mem_reg[33][40]  ( .D(n24803), .E(n6428), .CP(clk), .QN(n3810) );
  EDFD1 \Mem_reg[32][40]  ( .D(n24803), .E(n6427), .CP(clk), .QN(n3762) );
  EDFD1 \Mem_reg[31][40]  ( .D(n24803), .E(n6426), .CP(clk), .QN(n3714) );
  EDFD1 \Mem_reg[30][40]  ( .D(n24803), .E(n6425), .CP(clk), .QN(n3666) );
  EDFD1 \Mem_reg[29][40]  ( .D(n24803), .E(n6424), .CP(clk), .QN(n3618) );
  EDFD1 \Mem_reg[28][40]  ( .D(n24803), .E(n6423), .CP(clk), .QN(n3570) );
  EDFD1 \Mem_reg[27][40]  ( .D(n24803), .E(n6422), .CP(clk), .QN(n3522) );
  EDFD1 \Mem_reg[26][40]  ( .D(n24803), .E(n6421), .CP(clk), .QN(n3474) );
  EDFD1 \Mem_reg[25][40]  ( .D(n24803), .E(n6420), .CP(clk), .QN(n3426) );
  EDFD1 \Mem_reg[24][40]  ( .D(n24803), .E(n6463), .CP(clk), .QN(n3378) );
  EDFD1 \Mem_reg[23][40]  ( .D(n24803), .E(n6464), .CP(clk), .QN(n3330) );
  EDFD1 \Mem_reg[22][40]  ( .D(n24803), .E(n6465), .CP(clk), .QN(n3282) );
  EDFD1 \Mem_reg[21][40]  ( .D(n24803), .E(n6466), .CP(clk), .QN(n3234) );
  EDFD1 \Mem_reg[20][40]  ( .D(n24803), .E(n6467), .CP(clk), .QN(n3186) );
  EDFD1 \Mem_reg[19][40]  ( .D(n24803), .E(n6468), .CP(clk), .QN(n3138) );
  EDFD1 \Mem_reg[18][40]  ( .D(n24803), .E(n6469), .CP(clk), .QN(n3090) );
  EDFD1 \Mem_reg[17][40]  ( .D(n24803), .E(n6470), .CP(clk), .QN(n3042) );
  EDFD1 \Mem_reg[16][40]  ( .D(n24803), .E(n6471), .CP(clk), .QN(n2994) );
  EDFD1 \Mem_reg[15][40]  ( .D(n24803), .E(n6472), .CP(clk), .QN(n2946) );
  EDFD1 \Mem_reg[14][40]  ( .D(n24803), .E(n24720), .CP(clk), .QN(n2898) );
  EDFD1 \Mem_reg[13][40]  ( .D(n24803), .E(n24709), .CP(clk), .QN(n2850) );
  EDFD1 \Mem_reg[12][40]  ( .D(n24803), .E(n24717), .CP(clk), .QN(n2802) );
  EDFD1 \Mem_reg[11][40]  ( .D(n24803), .E(n24707), .CP(clk), .QN(n2754) );
  EDFD1 \Mem_reg[10][40]  ( .D(n24803), .E(n6477), .CP(clk), .QN(n2706) );
  EDFD1 \Mem_reg[9][40]  ( .D(n24803), .E(n24708), .CP(clk), .QN(n2658) );
  EDFD1 \Mem_reg[8][40]  ( .D(n24803), .E(n15642), .CP(clk), .QN(n2610) );
  EDFD1 \Mem_reg[7][40]  ( .D(n24803), .E(n24718), .CP(clk), .QN(n2562) );
  EDFD1 \Mem_reg[6][40]  ( .D(n24803), .E(n24716), .CP(clk), .QN(n2514) );
  EDFD1 \Mem_reg[5][40]  ( .D(n24803), .E(n24719), .CP(clk), .QN(n2466) );
  EDFD1 \Mem_reg[4][40]  ( .D(n24803), .E(n24706), .CP(clk), .QN(n2418) );
  EDFD1 \Mem_reg[3][40]  ( .D(n24803), .E(n24721), .CP(clk), .QN(n2370) );
  EDFD1 \Mem_reg[2][40]  ( .D(n24803), .E(n6460), .CP(clk), .QN(n2322) );
  EDFD1 \Mem_reg[1][40]  ( .D(n24803), .E(n24703), .CP(clk), .QN(n2274) );
  EDFD1 \Mem_reg[0][40]  ( .D(n24803), .E(n24705), .CP(clk), .QN(n2226) );
  EDFD1 \Mem_reg[88][39]  ( .D(n24801), .E(n6419), .CP(clk), .Q(n27193) );
  EDFD1 \Mem_reg[87][39]  ( .D(n24801), .E(n6418), .CP(clk), .QN(n6307) );
  EDFD1 \Mem_reg[86][39]  ( .D(n24801), .E(n6417), .CP(clk), .QN(n24676) );
  EDFD1 \Mem_reg[85][39]  ( .D(n24801), .E(n6416), .CP(clk), .QN(n6211) );
  EDFD1 \Mem_reg[84][39]  ( .D(n24801), .E(n6415), .CP(clk), .QN(n6163) );
  EDFD1 \Mem_reg[83][39]  ( .D(n24801), .E(n6414), .CP(clk), .QN(n6115) );
  EDFD1 \Mem_reg[82][39]  ( .D(n24801), .E(n6413), .CP(clk), .QN(n6067) );
  EDFD1 \Mem_reg[81][39]  ( .D(n24801), .E(n6412), .CP(clk), .QN(n6019) );
  EDFD1 \Mem_reg[80][39]  ( .D(n24801), .E(n6411), .CP(clk), .QN(n5971) );
  EDFD1 \Mem_reg[79][39]  ( .D(n24801), .E(n6410), .CP(clk), .QN(n5923) );
  EDFD1 \Mem_reg[78][39]  ( .D(n24801), .E(n6409), .CP(clk), .QN(n5875) );
  EDFD1 \Mem_reg[77][39]  ( .D(n24801), .E(n6408), .CP(clk), .QN(n5827) );
  EDFD1 \Mem_reg[76][39]  ( .D(n24801), .E(n6407), .CP(clk), .QN(n5779) );
  EDFD1 \Mem_reg[75][39]  ( .D(n24801), .E(n6406), .CP(clk), .QN(n27194) );
  EDFD1 \Mem_reg[74][39]  ( .D(n24801), .E(n6405), .CP(clk), .QN(n5683) );
  EDFD1 \Mem_reg[73][39]  ( .D(n24801), .E(n6404), .CP(clk), .QN(n27195) );
  EDFD1 \Mem_reg[72][39]  ( .D(n24801), .E(n6403), .CP(clk), .QN(n5587) );
  EDFD1 \Mem_reg[71][39]  ( .D(n24801), .E(n6402), .CP(clk), .QN(n5539) );
  EDFD1 \Mem_reg[70][39]  ( .D(n24801), .E(n6401), .CP(clk), .QN(n5491) );
  EDFD1 \Mem_reg[69][39]  ( .D(n24801), .E(n6400), .CP(clk), .QN(n5443) );
  EDFD1 \Mem_reg[68][39]  ( .D(n24801), .E(n6399), .CP(clk), .QN(n5395) );
  EDFD1 \Mem_reg[67][39]  ( .D(n24801), .E(n6398), .CP(clk), .QN(n5347) );
  EDFD1 \Mem_reg[66][39]  ( .D(n24801), .E(n6397), .CP(clk), .QN(n5299) );
  EDFD1 \Mem_reg[65][39]  ( .D(n24801), .E(n6396), .CP(clk), .QN(n15605) );
  EDFD1 \Mem_reg[64][39]  ( .D(n24801), .E(n6395), .CP(clk), .QN(n5203) );
  EDFD1 \Mem_reg[63][39]  ( .D(n24801), .E(n6456), .CP(clk), .QN(n5155) );
  EDFD1 \Mem_reg[62][39]  ( .D(n24801), .E(n6455), .CP(clk), .QN(n5107) );
  EDFD1 \Mem_reg[61][39]  ( .D(n24801), .E(n6454), .CP(clk), .QN(n18044) );
  EDFD1 \Mem_reg[60][39]  ( .D(n24801), .E(n6453), .CP(clk), .QN(n18043) );
  EDFD1 \Mem_reg[59][39]  ( .D(n24801), .E(n6452), .CP(clk), .QN(n4963) );
  EDFD1 \Mem_reg[58][39]  ( .D(n24801), .E(n6451), .CP(clk), .QN(n4915) );
  EDFD1 \Mem_reg[57][39]  ( .D(n24801), .E(n6450), .CP(clk), .QN(n4867) );
  EDFD1 \Mem_reg[56][39]  ( .D(n24801), .E(n6449), .CP(clk), .QN(n4819) );
  EDFD1 \Mem_reg[55][39]  ( .D(n24801), .E(n6448), .CP(clk), .QN(n4771) );
  EDFD1 \Mem_reg[54][39]  ( .D(n24801), .E(n6447), .CP(clk), .QN(n15604) );
  EDFD1 \Mem_reg[53][39]  ( .D(n24801), .E(n6446), .CP(clk), .QN(n4675) );
  EDFD1 \Mem_reg[52][39]  ( .D(n24801), .E(n6445), .CP(clk), .Q(n27192) );
  EDFD1 \Mem_reg[51][39]  ( .D(n24801), .E(n6444), .CP(clk), .QN(n4579) );
  EDFD1 \Mem_reg[50][39]  ( .D(n24801), .E(n6443), .CP(clk), .QN(n4531) );
  EDFD1 \Mem_reg[49][39]  ( .D(n24801), .E(n6442), .CP(clk), .QN(n4483) );
  EDFD1 \Mem_reg[48][39]  ( .D(n24801), .E(n6441), .CP(clk), .QN(n4435) );
  EDFD1 \Mem_reg[47][39]  ( .D(n24801), .E(n6440), .CP(clk), .QN(n4387) );
  EDFD1 \Mem_reg[46][39]  ( .D(n24801), .E(n6439), .CP(clk), .QN(n4339) );
  EDFD1 \Mem_reg[43][39]  ( .D(n24801), .E(n6438), .CP(clk), .QN(n4291) );
  EDFD1 \Mem_reg[42][39]  ( .D(n24801), .E(n6437), .CP(clk), .QN(n4243) );
  EDFD1 \Mem_reg[41][39]  ( .D(n24801), .E(n6436), .CP(clk), .QN(n4195) );
  EDFD1 \Mem_reg[40][39]  ( .D(n24801), .E(n6435), .CP(clk), .QN(n4147) );
  EDFD1 \Mem_reg[39][39]  ( .D(n24801), .E(n6434), .CP(clk), .QN(n4099) );
  EDFD1 \Mem_reg[38][39]  ( .D(n24801), .E(n6433), .CP(clk), .QN(n4051) );
  EDFD1 \Mem_reg[37][39]  ( .D(n24801), .E(n6432), .CP(clk), .QN(n4003) );
  EDFD1 \Mem_reg[36][39]  ( .D(n24801), .E(n6431), .CP(clk), .QN(n3955) );
  EDFD1 \Mem_reg[35][39]  ( .D(n24801), .E(n6430), .CP(clk), .QN(n3907) );
  EDFD1 \Mem_reg[34][39]  ( .D(n24801), .E(n6429), .CP(clk), .QN(n3859) );
  EDFD1 \Mem_reg[33][39]  ( .D(n24801), .E(n6428), .CP(clk), .QN(n3811) );
  EDFD1 \Mem_reg[32][39]  ( .D(n24801), .E(n6427), .CP(clk), .QN(n3763) );
  EDFD1 \Mem_reg[31][39]  ( .D(n24801), .E(n6426), .CP(clk), .QN(n3715) );
  EDFD1 \Mem_reg[30][39]  ( .D(n24801), .E(n6425), .CP(clk), .QN(n3667) );
  EDFD1 \Mem_reg[29][39]  ( .D(n24801), .E(n6424), .CP(clk), .QN(n3619) );
  EDFD1 \Mem_reg[28][39]  ( .D(n24801), .E(n6423), .CP(clk), .QN(n3571) );
  EDFD1 \Mem_reg[27][39]  ( .D(n24801), .E(n6422), .CP(clk), .QN(n3523) );
  EDFD1 \Mem_reg[26][39]  ( .D(n24801), .E(n6421), .CP(clk), .QN(n3475) );
  EDFD1 \Mem_reg[25][39]  ( .D(n24801), .E(n6420), .CP(clk), .QN(n3427) );
  EDFD1 \Mem_reg[24][39]  ( .D(n24801), .E(n6463), .CP(clk), .QN(n3379) );
  EDFD1 \Mem_reg[23][39]  ( .D(n24801), .E(n6464), .CP(clk), .QN(n3331) );
  EDFD1 \Mem_reg[22][39]  ( .D(n24801), .E(n6465), .CP(clk), .QN(n3283) );
  EDFD1 \Mem_reg[21][39]  ( .D(n24801), .E(n6466), .CP(clk), .QN(n3235) );
  EDFD1 \Mem_reg[20][39]  ( .D(n24801), .E(n6467), .CP(clk), .QN(n3187) );
  EDFD1 \Mem_reg[19][39]  ( .D(n24801), .E(n6468), .CP(clk), .QN(n3139) );
  EDFD1 \Mem_reg[18][39]  ( .D(n24801), .E(n6469), .CP(clk), .QN(n3091) );
  EDFD1 \Mem_reg[17][39]  ( .D(n24801), .E(n6470), .CP(clk), .QN(n3043) );
  EDFD1 \Mem_reg[16][39]  ( .D(n24801), .E(n6471), .CP(clk), .QN(n2995) );
  EDFD1 \Mem_reg[15][39]  ( .D(n24801), .E(n6472), .CP(clk), .QN(n2947) );
  EDFD1 \Mem_reg[14][39]  ( .D(n24801), .E(n24720), .CP(clk), .QN(n2899) );
  EDFD1 \Mem_reg[13][39]  ( .D(n24801), .E(n24709), .CP(clk), .QN(n2851) );
  EDFD1 \Mem_reg[12][39]  ( .D(n24801), .E(n24717), .CP(clk), .QN(n2803) );
  EDFD1 \Mem_reg[11][39]  ( .D(n24801), .E(n24707), .CP(clk), .QN(n2755) );
  EDFD1 \Mem_reg[10][39]  ( .D(n24801), .E(n6477), .CP(clk), .QN(n2707) );
  EDFD1 \Mem_reg[9][39]  ( .D(n24801), .E(n24708), .CP(clk), .QN(n2659) );
  EDFD1 \Mem_reg[8][39]  ( .D(n24801), .E(n15642), .CP(clk), .QN(n2611) );
  EDFD1 \Mem_reg[7][39]  ( .D(n24801), .E(n24718), .CP(clk), .QN(n2563) );
  EDFD1 \Mem_reg[6][39]  ( .D(n24801), .E(n24716), .CP(clk), .QN(n2515) );
  EDFD1 \Mem_reg[5][39]  ( .D(n24801), .E(n24719), .CP(clk), .QN(n2467) );
  EDFD1 \Mem_reg[4][39]  ( .D(n24801), .E(n24706), .CP(clk), .QN(n2419) );
  EDFD1 \Mem_reg[3][39]  ( .D(n24801), .E(n24721), .CP(clk), .QN(n2371) );
  EDFD1 \Mem_reg[2][39]  ( .D(n24801), .E(n6460), .CP(clk), .QN(n2323) );
  EDFD1 \Mem_reg[1][39]  ( .D(n24801), .E(n24703), .CP(clk), .QN(n2275) );
  EDFD1 \Mem_reg[0][39]  ( .D(n24801), .E(n24705), .CP(clk), .QN(n2227) );
  EDFD1 \Mem_reg[88][38]  ( .D(n24799), .E(n6419), .CP(clk), .Q(n27189) );
  EDFD1 \Mem_reg[87][38]  ( .D(n24799), .E(n6418), .CP(clk), .QN(n6308) );
  EDFD1 \Mem_reg[86][38]  ( .D(n24799), .E(n6417), .CP(clk), .QN(n24673) );
  EDFD1 \Mem_reg[85][38]  ( .D(n24799), .E(n6416), .CP(clk), .QN(n6212) );
  EDFD1 \Mem_reg[84][38]  ( .D(n24799), .E(n6415), .CP(clk), .QN(n6164) );
  EDFD1 \Mem_reg[83][38]  ( .D(n24799), .E(n6414), .CP(clk), .QN(n6116) );
  EDFD1 \Mem_reg[82][38]  ( .D(n24799), .E(n6413), .CP(clk), .QN(n6068) );
  EDFD1 \Mem_reg[81][38]  ( .D(n24799), .E(n6412), .CP(clk), .QN(n6020) );
  EDFD1 \Mem_reg[80][38]  ( .D(n24799), .E(n6411), .CP(clk), .QN(n5972) );
  EDFD1 \Mem_reg[79][38]  ( .D(n24799), .E(n6410), .CP(clk), .QN(n5924) );
  EDFD1 \Mem_reg[78][38]  ( .D(n24799), .E(n6409), .CP(clk), .QN(n5876) );
  EDFD1 \Mem_reg[77][38]  ( .D(n24799), .E(n6408), .CP(clk), .QN(n5828) );
  EDFD1 \Mem_reg[76][38]  ( .D(n24799), .E(n6407), .CP(clk), .QN(n5780) );
  EDFD1 \Mem_reg[75][38]  ( .D(n24799), .E(n6406), .CP(clk), .QN(n27190) );
  EDFD1 \Mem_reg[74][38]  ( .D(n24799), .E(n6405), .CP(clk), .QN(n5684) );
  EDFD1 \Mem_reg[73][38]  ( .D(n24799), .E(n6404), .CP(clk), .QN(n27191) );
  EDFD1 \Mem_reg[72][38]  ( .D(n24799), .E(n6403), .CP(clk), .QN(n5588) );
  EDFD1 \Mem_reg[71][38]  ( .D(n24799), .E(n6402), .CP(clk), .QN(n5540) );
  EDFD1 \Mem_reg[70][38]  ( .D(n24799), .E(n6401), .CP(clk), .QN(n5492) );
  EDFD1 \Mem_reg[69][38]  ( .D(n24799), .E(n6400), .CP(clk), .QN(n5444) );
  EDFD1 \Mem_reg[68][38]  ( .D(n24799), .E(n6399), .CP(clk), .QN(n5396) );
  EDFD1 \Mem_reg[67][38]  ( .D(n24799), .E(n6398), .CP(clk), .QN(n5348) );
  EDFD1 \Mem_reg[66][38]  ( .D(n24799), .E(n6397), .CP(clk), .QN(n5300) );
  EDFD1 \Mem_reg[65][38]  ( .D(n24799), .E(n6396), .CP(clk), .QN(n15601) );
  EDFD1 \Mem_reg[64][38]  ( .D(n24799), .E(n6395), .CP(clk), .QN(n5204) );
  EDFD1 \Mem_reg[63][38]  ( .D(n24799), .E(n6456), .CP(clk), .QN(n5156) );
  EDFD1 \Mem_reg[62][38]  ( .D(n24799), .E(n6455), .CP(clk), .QN(n5108) );
  EDFD1 \Mem_reg[61][38]  ( .D(n24799), .E(n6454), .CP(clk), .QN(n18041) );
  EDFD1 \Mem_reg[60][38]  ( .D(n24799), .E(n6453), .CP(clk), .QN(n18040) );
  EDFD1 \Mem_reg[59][38]  ( .D(n24799), .E(n6452), .CP(clk), .QN(n4964) );
  EDFD1 \Mem_reg[58][38]  ( .D(n24799), .E(n6451), .CP(clk), .QN(n4916) );
  EDFD1 \Mem_reg[57][38]  ( .D(n24799), .E(n6450), .CP(clk), .QN(n4868) );
  EDFD1 \Mem_reg[56][38]  ( .D(n24799), .E(n6449), .CP(clk), .QN(n4820) );
  EDFD1 \Mem_reg[55][38]  ( .D(n24799), .E(n6448), .CP(clk), .QN(n4772) );
  EDFD1 \Mem_reg[54][38]  ( .D(n24799), .E(n6447), .CP(clk), .QN(n15600) );
  EDFD1 \Mem_reg[53][38]  ( .D(n24799), .E(n6446), .CP(clk), .QN(n4676) );
  EDFD1 \Mem_reg[52][38]  ( .D(n24799), .E(n6445), .CP(clk), .Q(n27188) );
  EDFD1 \Mem_reg[51][38]  ( .D(n24799), .E(n6444), .CP(clk), .QN(n4580) );
  EDFD1 \Mem_reg[50][38]  ( .D(n24799), .E(n6443), .CP(clk), .QN(n4532) );
  EDFD1 \Mem_reg[49][38]  ( .D(n24799), .E(n6442), .CP(clk), .QN(n4484) );
  EDFD1 \Mem_reg[48][38]  ( .D(n24799), .E(n6441), .CP(clk), .QN(n4436) );
  EDFD1 \Mem_reg[47][38]  ( .D(n24799), .E(n6440), .CP(clk), .QN(n4388) );
  EDFD1 \Mem_reg[46][38]  ( .D(n24799), .E(n6439), .CP(clk), .QN(n4340) );
  EDFD1 \Mem_reg[43][38]  ( .D(n24799), .E(n6438), .CP(clk), .QN(n4292) );
  EDFD1 \Mem_reg[42][38]  ( .D(n24799), .E(n6437), .CP(clk), .QN(n4244) );
  EDFD1 \Mem_reg[41][38]  ( .D(n24799), .E(n6436), .CP(clk), .QN(n4196) );
  EDFD1 \Mem_reg[40][38]  ( .D(n24799), .E(n6435), .CP(clk), .QN(n4148) );
  EDFD1 \Mem_reg[39][38]  ( .D(n24799), .E(n6434), .CP(clk), .QN(n4100) );
  EDFD1 \Mem_reg[38][38]  ( .D(n24799), .E(n6433), .CP(clk), .QN(n4052) );
  EDFD1 \Mem_reg[37][38]  ( .D(n24799), .E(n6432), .CP(clk), .QN(n4004) );
  EDFD1 \Mem_reg[36][38]  ( .D(n24799), .E(n6431), .CP(clk), .QN(n3956) );
  EDFD1 \Mem_reg[35][38]  ( .D(n24799), .E(n6430), .CP(clk), .QN(n3908) );
  EDFD1 \Mem_reg[34][38]  ( .D(n24799), .E(n6429), .CP(clk), .QN(n3860) );
  EDFD1 \Mem_reg[33][38]  ( .D(n24799), .E(n6428), .CP(clk), .QN(n3812) );
  EDFD1 \Mem_reg[32][38]  ( .D(n24799), .E(n6427), .CP(clk), .QN(n3764) );
  EDFD1 \Mem_reg[31][38]  ( .D(n24799), .E(n6426), .CP(clk), .QN(n3716) );
  EDFD1 \Mem_reg[30][38]  ( .D(n24799), .E(n6425), .CP(clk), .QN(n3668) );
  EDFD1 \Mem_reg[29][38]  ( .D(n24799), .E(n6424), .CP(clk), .QN(n3620) );
  EDFD1 \Mem_reg[28][38]  ( .D(n24799), .E(n6423), .CP(clk), .QN(n3572) );
  EDFD1 \Mem_reg[27][38]  ( .D(n24799), .E(n6422), .CP(clk), .QN(n3524) );
  EDFD1 \Mem_reg[26][38]  ( .D(n24799), .E(n6421), .CP(clk), .QN(n3476) );
  EDFD1 \Mem_reg[25][38]  ( .D(n24799), .E(n6420), .CP(clk), .QN(n3428) );
  EDFD1 \Mem_reg[24][38]  ( .D(n24799), .E(n6463), .CP(clk), .QN(n3380) );
  EDFD1 \Mem_reg[23][38]  ( .D(n24799), .E(n6464), .CP(clk), .QN(n3332) );
  EDFD1 \Mem_reg[22][38]  ( .D(n24799), .E(n6465), .CP(clk), .QN(n3284) );
  EDFD1 \Mem_reg[21][38]  ( .D(n24799), .E(n6466), .CP(clk), .QN(n3236) );
  EDFD1 \Mem_reg[20][38]  ( .D(n24799), .E(n6467), .CP(clk), .QN(n3188) );
  EDFD1 \Mem_reg[19][38]  ( .D(n24799), .E(n6468), .CP(clk), .QN(n3140) );
  EDFD1 \Mem_reg[18][38]  ( .D(n24799), .E(n6469), .CP(clk), .QN(n3092) );
  EDFD1 \Mem_reg[17][38]  ( .D(n24799), .E(n6470), .CP(clk), .QN(n3044) );
  EDFD1 \Mem_reg[16][38]  ( .D(n24799), .E(n6471), .CP(clk), .QN(n2996) );
  EDFD1 \Mem_reg[15][38]  ( .D(n24799), .E(n6472), .CP(clk), .QN(n2948) );
  EDFD1 \Mem_reg[14][38]  ( .D(n24799), .E(n24720), .CP(clk), .QN(n2900) );
  EDFD1 \Mem_reg[13][38]  ( .D(n24799), .E(n24709), .CP(clk), .QN(n2852) );
  EDFD1 \Mem_reg[12][38]  ( .D(n24799), .E(n24717), .CP(clk), .QN(n2804) );
  EDFD1 \Mem_reg[11][38]  ( .D(n24799), .E(n24707), .CP(clk), .QN(n2756) );
  EDFD1 \Mem_reg[10][38]  ( .D(n24799), .E(n6477), .CP(clk), .QN(n2708) );
  EDFD1 \Mem_reg[9][38]  ( .D(n24799), .E(n24708), .CP(clk), .QN(n2660) );
  EDFD1 \Mem_reg[8][38]  ( .D(n24799), .E(n15642), .CP(clk), .QN(n2612) );
  EDFD1 \Mem_reg[7][38]  ( .D(n24799), .E(n24718), .CP(clk), .QN(n2564) );
  EDFD1 \Mem_reg[6][38]  ( .D(n24799), .E(n24716), .CP(clk), .QN(n2516) );
  EDFD1 \Mem_reg[5][38]  ( .D(n24799), .E(n24719), .CP(clk), .QN(n2468) );
  EDFD1 \Mem_reg[4][38]  ( .D(n24799), .E(n24706), .CP(clk), .QN(n2420) );
  EDFD1 \Mem_reg[3][38]  ( .D(n24799), .E(n24721), .CP(clk), .QN(n2372) );
  EDFD1 \Mem_reg[2][38]  ( .D(n24799), .E(n6460), .CP(clk), .QN(n2324) );
  EDFD1 \Mem_reg[1][38]  ( .D(n24799), .E(n24703), .CP(clk), .QN(n2276) );
  EDFD1 \Mem_reg[0][38]  ( .D(n24799), .E(n24705), .CP(clk), .QN(n2228) );
  EDFD1 \Mem_reg[88][37]  ( .D(n24797), .E(n6419), .CP(clk), .Q(n27185) );
  EDFD1 \Mem_reg[87][37]  ( .D(n24797), .E(n6418), .CP(clk), .QN(n6309) );
  EDFD1 \Mem_reg[86][37]  ( .D(n24797), .E(n6417), .CP(clk), .QN(n24670) );
  EDFD1 \Mem_reg[85][37]  ( .D(n24797), .E(n6416), .CP(clk), .QN(n6213) );
  EDFD1 \Mem_reg[84][37]  ( .D(n24797), .E(n6415), .CP(clk), .QN(n6165) );
  EDFD1 \Mem_reg[83][37]  ( .D(n24797), .E(n6414), .CP(clk), .QN(n6117) );
  EDFD1 \Mem_reg[82][37]  ( .D(n24797), .E(n6413), .CP(clk), .QN(n6069) );
  EDFD1 \Mem_reg[81][37]  ( .D(n24797), .E(n6412), .CP(clk), .QN(n6021) );
  EDFD1 \Mem_reg[80][37]  ( .D(n24797), .E(n6411), .CP(clk), .QN(n5973) );
  EDFD1 \Mem_reg[79][37]  ( .D(n24797), .E(n6410), .CP(clk), .QN(n5925) );
  EDFD1 \Mem_reg[78][37]  ( .D(n24797), .E(n6409), .CP(clk), .QN(n5877) );
  EDFD1 \Mem_reg[77][37]  ( .D(n24797), .E(n6408), .CP(clk), .QN(n5829) );
  EDFD1 \Mem_reg[76][37]  ( .D(n24797), .E(n6407), .CP(clk), .QN(n5781) );
  EDFD1 \Mem_reg[75][37]  ( .D(n24797), .E(n6406), .CP(clk), .QN(n27186) );
  EDFD1 \Mem_reg[74][37]  ( .D(n24797), .E(n6405), .CP(clk), .QN(n5685) );
  EDFD1 \Mem_reg[73][37]  ( .D(n24797), .E(n6404), .CP(clk), .QN(n27187) );
  EDFD1 \Mem_reg[72][37]  ( .D(n24797), .E(n6403), .CP(clk), .QN(n5589) );
  EDFD1 \Mem_reg[71][37]  ( .D(n24797), .E(n6402), .CP(clk), .QN(n5541) );
  EDFD1 \Mem_reg[70][37]  ( .D(n24797), .E(n6401), .CP(clk), .QN(n5493) );
  EDFD1 \Mem_reg[69][37]  ( .D(n24797), .E(n6400), .CP(clk), .QN(n5445) );
  EDFD1 \Mem_reg[68][37]  ( .D(n24797), .E(n6399), .CP(clk), .QN(n5397) );
  EDFD1 \Mem_reg[67][37]  ( .D(n24797), .E(n6398), .CP(clk), .QN(n5349) );
  EDFD1 \Mem_reg[66][37]  ( .D(n24797), .E(n6397), .CP(clk), .QN(n5301) );
  EDFD1 \Mem_reg[65][37]  ( .D(n24797), .E(n6396), .CP(clk), .QN(n15597) );
  EDFD1 \Mem_reg[64][37]  ( .D(n24797), .E(n6395), .CP(clk), .QN(n5205) );
  EDFD1 \Mem_reg[63][37]  ( .D(n24797), .E(n6456), .CP(clk), .QN(n5157) );
  EDFD1 \Mem_reg[62][37]  ( .D(n24797), .E(n6455), .CP(clk), .QN(n5109) );
  EDFD1 \Mem_reg[61][37]  ( .D(n24797), .E(n6454), .CP(clk), .QN(n18038) );
  EDFD1 \Mem_reg[60][37]  ( .D(n24797), .E(n6453), .CP(clk), .QN(n18037) );
  EDFD1 \Mem_reg[59][37]  ( .D(n24797), .E(n6452), .CP(clk), .QN(n4965) );
  EDFD1 \Mem_reg[58][37]  ( .D(n24797), .E(n6451), .CP(clk), .QN(n4917) );
  EDFD1 \Mem_reg[57][37]  ( .D(n24797), .E(n6450), .CP(clk), .QN(n4869) );
  EDFD1 \Mem_reg[56][37]  ( .D(n24797), .E(n6449), .CP(clk), .QN(n4821) );
  EDFD1 \Mem_reg[55][37]  ( .D(n24797), .E(n6448), .CP(clk), .QN(n4773) );
  EDFD1 \Mem_reg[54][37]  ( .D(n24797), .E(n6447), .CP(clk), .QN(n15596) );
  EDFD1 \Mem_reg[53][37]  ( .D(n24797), .E(n6446), .CP(clk), .QN(n4677) );
  EDFD1 \Mem_reg[52][37]  ( .D(n24797), .E(n6445), .CP(clk), .Q(n27184) );
  EDFD1 \Mem_reg[51][37]  ( .D(n24797), .E(n6444), .CP(clk), .QN(n4581) );
  EDFD1 \Mem_reg[50][37]  ( .D(n24797), .E(n6443), .CP(clk), .QN(n4533) );
  EDFD1 \Mem_reg[49][37]  ( .D(n24797), .E(n6442), .CP(clk), .QN(n4485) );
  EDFD1 \Mem_reg[48][37]  ( .D(n24797), .E(n6441), .CP(clk), .QN(n4437) );
  EDFD1 \Mem_reg[47][37]  ( .D(n24797), .E(n6440), .CP(clk), .QN(n4389) );
  EDFD1 \Mem_reg[46][37]  ( .D(n24797), .E(n6439), .CP(clk), .QN(n4341) );
  EDFD1 \Mem_reg[43][37]  ( .D(n24797), .E(n6438), .CP(clk), .QN(n4293) );
  EDFD1 \Mem_reg[42][37]  ( .D(n24797), .E(n6437), .CP(clk), .QN(n4245) );
  EDFD1 \Mem_reg[41][37]  ( .D(n24797), .E(n6436), .CP(clk), .QN(n4197) );
  EDFD1 \Mem_reg[40][37]  ( .D(n24797), .E(n6435), .CP(clk), .QN(n4149) );
  EDFD1 \Mem_reg[39][37]  ( .D(n24797), .E(n6434), .CP(clk), .QN(n4101) );
  EDFD1 \Mem_reg[38][37]  ( .D(n24797), .E(n6433), .CP(clk), .QN(n4053) );
  EDFD1 \Mem_reg[37][37]  ( .D(n24797), .E(n6432), .CP(clk), .QN(n4005) );
  EDFD1 \Mem_reg[36][37]  ( .D(n24797), .E(n6431), .CP(clk), .QN(n3957) );
  EDFD1 \Mem_reg[35][37]  ( .D(n24797), .E(n6430), .CP(clk), .QN(n3909) );
  EDFD1 \Mem_reg[34][37]  ( .D(n24797), .E(n6429), .CP(clk), .QN(n3861) );
  EDFD1 \Mem_reg[33][37]  ( .D(n24797), .E(n6428), .CP(clk), .QN(n3813) );
  EDFD1 \Mem_reg[32][37]  ( .D(n24797), .E(n6427), .CP(clk), .QN(n3765) );
  EDFD1 \Mem_reg[31][37]  ( .D(n24797), .E(n6426), .CP(clk), .QN(n3717) );
  EDFD1 \Mem_reg[30][37]  ( .D(n24797), .E(n6425), .CP(clk), .QN(n3669) );
  EDFD1 \Mem_reg[29][37]  ( .D(n24797), .E(n6424), .CP(clk), .QN(n3621) );
  EDFD1 \Mem_reg[28][37]  ( .D(n24797), .E(n6423), .CP(clk), .QN(n3573) );
  EDFD1 \Mem_reg[27][37]  ( .D(n24797), .E(n6422), .CP(clk), .QN(n3525) );
  EDFD1 \Mem_reg[26][37]  ( .D(n24797), .E(n6421), .CP(clk), .QN(n3477) );
  EDFD1 \Mem_reg[25][37]  ( .D(n24797), .E(n6420), .CP(clk), .QN(n3429) );
  EDFD1 \Mem_reg[24][37]  ( .D(n24797), .E(n6463), .CP(clk), .QN(n3381) );
  EDFD1 \Mem_reg[23][37]  ( .D(n24797), .E(n6464), .CP(clk), .QN(n3333) );
  EDFD1 \Mem_reg[22][37]  ( .D(n24797), .E(n6465), .CP(clk), .QN(n3285) );
  EDFD1 \Mem_reg[21][37]  ( .D(n24797), .E(n6466), .CP(clk), .QN(n3237) );
  EDFD1 \Mem_reg[20][37]  ( .D(n24797), .E(n6467), .CP(clk), .QN(n3189) );
  EDFD1 \Mem_reg[19][37]  ( .D(n24797), .E(n6468), .CP(clk), .QN(n3141) );
  EDFD1 \Mem_reg[18][37]  ( .D(n24797), .E(n6469), .CP(clk), .QN(n3093) );
  EDFD1 \Mem_reg[17][37]  ( .D(n24797), .E(n6470), .CP(clk), .QN(n3045) );
  EDFD1 \Mem_reg[16][37]  ( .D(n24797), .E(n6471), .CP(clk), .QN(n2997) );
  EDFD1 \Mem_reg[15][37]  ( .D(n24797), .E(n6472), .CP(clk), .QN(n2949) );
  EDFD1 \Mem_reg[14][37]  ( .D(n24797), .E(n24720), .CP(clk), .QN(n2901) );
  EDFD1 \Mem_reg[13][37]  ( .D(n24797), .E(n24709), .CP(clk), .QN(n2853) );
  EDFD1 \Mem_reg[12][37]  ( .D(n24797), .E(n24717), .CP(clk), .QN(n2805) );
  EDFD1 \Mem_reg[11][37]  ( .D(n24797), .E(n24707), .CP(clk), .QN(n2757) );
  EDFD1 \Mem_reg[10][37]  ( .D(n24797), .E(n6477), .CP(clk), .QN(n2709) );
  EDFD1 \Mem_reg[9][37]  ( .D(n24797), .E(n24708), .CP(clk), .QN(n2661) );
  EDFD1 \Mem_reg[8][37]  ( .D(n24797), .E(n15642), .CP(clk), .QN(n2613) );
  EDFD1 \Mem_reg[7][37]  ( .D(n24797), .E(n24718), .CP(clk), .QN(n2565) );
  EDFD1 \Mem_reg[6][37]  ( .D(n24797), .E(n24716), .CP(clk), .QN(n2517) );
  EDFD1 \Mem_reg[5][37]  ( .D(n24797), .E(n24719), .CP(clk), .QN(n2469) );
  EDFD1 \Mem_reg[4][37]  ( .D(n24797), .E(n24706), .CP(clk), .QN(n2421) );
  EDFD1 \Mem_reg[3][37]  ( .D(n24797), .E(n24721), .CP(clk), .QN(n2373) );
  EDFD1 \Mem_reg[2][37]  ( .D(n24797), .E(n6460), .CP(clk), .QN(n2325) );
  EDFD1 \Mem_reg[1][37]  ( .D(n24797), .E(n24703), .CP(clk), .QN(n2277) );
  EDFD1 \Mem_reg[0][37]  ( .D(n24797), .E(n24705), .CP(clk), .QN(n2229) );
  EDFD1 \Mem_reg[88][36]  ( .D(n24795), .E(n6419), .CP(clk), .Q(n27181) );
  EDFD1 \Mem_reg[87][36]  ( .D(n24795), .E(n6418), .CP(clk), .QN(n6310) );
  EDFD1 \Mem_reg[86][36]  ( .D(n24795), .E(n6417), .CP(clk), .QN(n24667) );
  EDFD1 \Mem_reg[85][36]  ( .D(n24795), .E(n6416), .CP(clk), .QN(n6214) );
  EDFD1 \Mem_reg[84][36]  ( .D(n24795), .E(n6415), .CP(clk), .QN(n6166) );
  EDFD1 \Mem_reg[83][36]  ( .D(n24795), .E(n6414), .CP(clk), .QN(n6118) );
  EDFD1 \Mem_reg[82][36]  ( .D(n24795), .E(n6413), .CP(clk), .QN(n6070) );
  EDFD1 \Mem_reg[81][36]  ( .D(n24795), .E(n6412), .CP(clk), .QN(n6022) );
  EDFD1 \Mem_reg[80][36]  ( .D(n24795), .E(n6411), .CP(clk), .QN(n5974) );
  EDFD1 \Mem_reg[79][36]  ( .D(n24795), .E(n6410), .CP(clk), .QN(n5926) );
  EDFD1 \Mem_reg[78][36]  ( .D(n24795), .E(n6409), .CP(clk), .QN(n5878) );
  EDFD1 \Mem_reg[77][36]  ( .D(n24795), .E(n6408), .CP(clk), .QN(n5830) );
  EDFD1 \Mem_reg[76][36]  ( .D(n24795), .E(n6407), .CP(clk), .QN(n5782) );
  EDFD1 \Mem_reg[75][36]  ( .D(n24795), .E(n6406), .CP(clk), .QN(n27182) );
  EDFD1 \Mem_reg[74][36]  ( .D(n24795), .E(n6405), .CP(clk), .QN(n5686) );
  EDFD1 \Mem_reg[73][36]  ( .D(n24795), .E(n6404), .CP(clk), .QN(n27183) );
  EDFD1 \Mem_reg[72][36]  ( .D(n24795), .E(n6403), .CP(clk), .QN(n5590) );
  EDFD1 \Mem_reg[71][36]  ( .D(n24795), .E(n6402), .CP(clk), .QN(n5542) );
  EDFD1 \Mem_reg[70][36]  ( .D(n24795), .E(n6401), .CP(clk), .QN(n5494) );
  EDFD1 \Mem_reg[69][36]  ( .D(n24795), .E(n6400), .CP(clk), .QN(n5446) );
  EDFD1 \Mem_reg[68][36]  ( .D(n24795), .E(n6399), .CP(clk), .QN(n5398) );
  EDFD1 \Mem_reg[67][36]  ( .D(n24795), .E(n6398), .CP(clk), .QN(n5350) );
  EDFD1 \Mem_reg[66][36]  ( .D(n24795), .E(n6397), .CP(clk), .QN(n5302) );
  EDFD1 \Mem_reg[65][36]  ( .D(n24795), .E(n6396), .CP(clk), .QN(n15593) );
  EDFD1 \Mem_reg[64][36]  ( .D(n24795), .E(n6395), .CP(clk), .QN(n5206) );
  EDFD1 \Mem_reg[63][36]  ( .D(n24795), .E(n6456), .CP(clk), .QN(n5158) );
  EDFD1 \Mem_reg[62][36]  ( .D(n24795), .E(n6455), .CP(clk), .QN(n5110) );
  EDFD1 \Mem_reg[61][36]  ( .D(n24795), .E(n6454), .CP(clk), .QN(n18035) );
  EDFD1 \Mem_reg[60][36]  ( .D(n24795), .E(n6453), .CP(clk), .QN(n18034) );
  EDFD1 \Mem_reg[59][36]  ( .D(n24795), .E(n6452), .CP(clk), .QN(n4966) );
  EDFD1 \Mem_reg[58][36]  ( .D(n24795), .E(n6451), .CP(clk), .QN(n4918) );
  EDFD1 \Mem_reg[57][36]  ( .D(n24795), .E(n6450), .CP(clk), .QN(n4870) );
  EDFD1 \Mem_reg[56][36]  ( .D(n24795), .E(n6449), .CP(clk), .QN(n4822) );
  EDFD1 \Mem_reg[55][36]  ( .D(n24795), .E(n6448), .CP(clk), .QN(n4774) );
  EDFD1 \Mem_reg[54][36]  ( .D(n24795), .E(n6447), .CP(clk), .QN(n15592) );
  EDFD1 \Mem_reg[53][36]  ( .D(n24795), .E(n6446), .CP(clk), .QN(n4678) );
  EDFD1 \Mem_reg[52][36]  ( .D(n24795), .E(n6445), .CP(clk), .Q(n27180) );
  EDFD1 \Mem_reg[51][36]  ( .D(n24795), .E(n6444), .CP(clk), .QN(n4582) );
  EDFD1 \Mem_reg[50][36]  ( .D(n24795), .E(n6443), .CP(clk), .QN(n4534) );
  EDFD1 \Mem_reg[49][36]  ( .D(n24795), .E(n6442), .CP(clk), .QN(n4486) );
  EDFD1 \Mem_reg[48][36]  ( .D(n24795), .E(n6441), .CP(clk), .QN(n4438) );
  EDFD1 \Mem_reg[47][36]  ( .D(n24795), .E(n6440), .CP(clk), .QN(n4390) );
  EDFD1 \Mem_reg[46][36]  ( .D(n24795), .E(n6439), .CP(clk), .QN(n4342) );
  EDFD1 \Mem_reg[43][36]  ( .D(n24795), .E(n6438), .CP(clk), .QN(n4294) );
  EDFD1 \Mem_reg[42][36]  ( .D(n24795), .E(n6437), .CP(clk), .QN(n4246) );
  EDFD1 \Mem_reg[41][36]  ( .D(n24795), .E(n6436), .CP(clk), .QN(n4198) );
  EDFD1 \Mem_reg[40][36]  ( .D(n24795), .E(n6435), .CP(clk), .QN(n4150) );
  EDFD1 \Mem_reg[39][36]  ( .D(n24795), .E(n6434), .CP(clk), .QN(n4102) );
  EDFD1 \Mem_reg[38][36]  ( .D(n24795), .E(n6433), .CP(clk), .QN(n4054) );
  EDFD1 \Mem_reg[37][36]  ( .D(n24795), .E(n6432), .CP(clk), .QN(n4006) );
  EDFD1 \Mem_reg[36][36]  ( .D(n24795), .E(n6431), .CP(clk), .QN(n3958) );
  EDFD1 \Mem_reg[35][36]  ( .D(n24795), .E(n6430), .CP(clk), .QN(n3910) );
  EDFD1 \Mem_reg[34][36]  ( .D(n24795), .E(n6429), .CP(clk), .QN(n3862) );
  EDFD1 \Mem_reg[33][36]  ( .D(n24795), .E(n6428), .CP(clk), .QN(n3814) );
  EDFD1 \Mem_reg[32][36]  ( .D(n24795), .E(n6427), .CP(clk), .QN(n3766) );
  EDFD1 \Mem_reg[31][36]  ( .D(n24795), .E(n6426), .CP(clk), .QN(n3718) );
  EDFD1 \Mem_reg[30][36]  ( .D(n24795), .E(n6425), .CP(clk), .QN(n3670) );
  EDFD1 \Mem_reg[29][36]  ( .D(n24795), .E(n6424), .CP(clk), .QN(n3622) );
  EDFD1 \Mem_reg[28][36]  ( .D(n24795), .E(n6423), .CP(clk), .QN(n3574) );
  EDFD1 \Mem_reg[27][36]  ( .D(n24795), .E(n6422), .CP(clk), .QN(n3526) );
  EDFD1 \Mem_reg[26][36]  ( .D(n24795), .E(n6421), .CP(clk), .QN(n3478) );
  EDFD1 \Mem_reg[25][36]  ( .D(n24795), .E(n6420), .CP(clk), .QN(n3430) );
  EDFD1 \Mem_reg[24][36]  ( .D(n24795), .E(n6463), .CP(clk), .QN(n3382) );
  EDFD1 \Mem_reg[23][36]  ( .D(n24795), .E(n6464), .CP(clk), .QN(n3334) );
  EDFD1 \Mem_reg[22][36]  ( .D(n24795), .E(n6465), .CP(clk), .QN(n3286) );
  EDFD1 \Mem_reg[21][36]  ( .D(n24795), .E(n6466), .CP(clk), .QN(n3238) );
  EDFD1 \Mem_reg[20][36]  ( .D(n24795), .E(n6467), .CP(clk), .QN(n3190) );
  EDFD1 \Mem_reg[19][36]  ( .D(n24795), .E(n6468), .CP(clk), .QN(n3142) );
  EDFD1 \Mem_reg[18][36]  ( .D(n24795), .E(n6469), .CP(clk), .QN(n3094) );
  EDFD1 \Mem_reg[17][36]  ( .D(n24795), .E(n6470), .CP(clk), .QN(n3046) );
  EDFD1 \Mem_reg[16][36]  ( .D(n24795), .E(n6471), .CP(clk), .QN(n2998) );
  EDFD1 \Mem_reg[15][36]  ( .D(n24795), .E(n6472), .CP(clk), .QN(n2950) );
  EDFD1 \Mem_reg[14][36]  ( .D(n24795), .E(n24720), .CP(clk), .QN(n2902) );
  EDFD1 \Mem_reg[13][36]  ( .D(n24795), .E(n24709), .CP(clk), .QN(n2854) );
  EDFD1 \Mem_reg[12][36]  ( .D(n24795), .E(n24717), .CP(clk), .QN(n2806) );
  EDFD1 \Mem_reg[11][36]  ( .D(n24795), .E(n24707), .CP(clk), .QN(n2758) );
  EDFD1 \Mem_reg[10][36]  ( .D(n24795), .E(n6477), .CP(clk), .QN(n2710) );
  EDFD1 \Mem_reg[9][36]  ( .D(n24795), .E(n24708), .CP(clk), .QN(n2662) );
  EDFD1 \Mem_reg[8][36]  ( .D(n24795), .E(n15642), .CP(clk), .QN(n2614) );
  EDFD1 \Mem_reg[7][36]  ( .D(n24795), .E(n24718), .CP(clk), .QN(n2566) );
  EDFD1 \Mem_reg[6][36]  ( .D(n24795), .E(n24716), .CP(clk), .QN(n2518) );
  EDFD1 \Mem_reg[5][36]  ( .D(n24795), .E(n24719), .CP(clk), .QN(n2470) );
  EDFD1 \Mem_reg[4][36]  ( .D(n24795), .E(n24706), .CP(clk), .QN(n2422) );
  EDFD1 \Mem_reg[3][36]  ( .D(n24795), .E(n24721), .CP(clk), .QN(n2374) );
  EDFD1 \Mem_reg[2][36]  ( .D(n24795), .E(n6460), .CP(clk), .QN(n2326) );
  EDFD1 \Mem_reg[1][36]  ( .D(n24795), .E(n24703), .CP(clk), .QN(n2278) );
  EDFD1 \Mem_reg[0][36]  ( .D(n24795), .E(n24705), .CP(clk), .QN(n2230) );
  EDFD1 \Mem_reg[88][35]  ( .D(n24793), .E(n6419), .CP(clk), .Q(n27177) );
  EDFD1 \Mem_reg[87][35]  ( .D(n24793), .E(n6418), .CP(clk), .QN(n6311) );
  EDFD1 \Mem_reg[86][35]  ( .D(n24793), .E(n6417), .CP(clk), .QN(n24664) );
  EDFD1 \Mem_reg[85][35]  ( .D(n24793), .E(n6416), .CP(clk), .QN(n6215) );
  EDFD1 \Mem_reg[84][35]  ( .D(n24793), .E(n6415), .CP(clk), .QN(n6167) );
  EDFD1 \Mem_reg[83][35]  ( .D(n24793), .E(n6414), .CP(clk), .QN(n6119) );
  EDFD1 \Mem_reg[82][35]  ( .D(n24793), .E(n6413), .CP(clk), .QN(n6071) );
  EDFD1 \Mem_reg[81][35]  ( .D(n24793), .E(n6412), .CP(clk), .QN(n6023) );
  EDFD1 \Mem_reg[80][35]  ( .D(n24793), .E(n6411), .CP(clk), .QN(n5975) );
  EDFD1 \Mem_reg[79][35]  ( .D(n24793), .E(n6410), .CP(clk), .QN(n5927) );
  EDFD1 \Mem_reg[78][35]  ( .D(n24793), .E(n6409), .CP(clk), .QN(n5879) );
  EDFD1 \Mem_reg[77][35]  ( .D(n24793), .E(n6408), .CP(clk), .QN(n5831) );
  EDFD1 \Mem_reg[76][35]  ( .D(n24793), .E(n6407), .CP(clk), .QN(n5783) );
  EDFD1 \Mem_reg[75][35]  ( .D(n24793), .E(n6406), .CP(clk), .QN(n27178) );
  EDFD1 \Mem_reg[74][35]  ( .D(n24793), .E(n6405), .CP(clk), .QN(n5687) );
  EDFD1 \Mem_reg[73][35]  ( .D(n24793), .E(n6404), .CP(clk), .QN(n27179) );
  EDFD1 \Mem_reg[72][35]  ( .D(n24793), .E(n6403), .CP(clk), .QN(n5591) );
  EDFD1 \Mem_reg[71][35]  ( .D(n24793), .E(n6402), .CP(clk), .QN(n5543) );
  EDFD1 \Mem_reg[70][35]  ( .D(n24793), .E(n6401), .CP(clk), .QN(n5495) );
  EDFD1 \Mem_reg[69][35]  ( .D(n24793), .E(n6400), .CP(clk), .QN(n5447) );
  EDFD1 \Mem_reg[68][35]  ( .D(n24793), .E(n6399), .CP(clk), .QN(n5399) );
  EDFD1 \Mem_reg[67][35]  ( .D(n24793), .E(n6398), .CP(clk), .QN(n5351) );
  EDFD1 \Mem_reg[66][35]  ( .D(n24793), .E(n6397), .CP(clk), .QN(n5303) );
  EDFD1 \Mem_reg[65][35]  ( .D(n24793), .E(n6396), .CP(clk), .QN(n15589) );
  EDFD1 \Mem_reg[64][35]  ( .D(n24793), .E(n6395), .CP(clk), .QN(n5207) );
  EDFD1 \Mem_reg[63][35]  ( .D(n24793), .E(n6456), .CP(clk), .QN(n5159) );
  EDFD1 \Mem_reg[62][35]  ( .D(n24793), .E(n6455), .CP(clk), .QN(n5111) );
  EDFD1 \Mem_reg[61][35]  ( .D(n24793), .E(n6454), .CP(clk), .QN(n18032) );
  EDFD1 \Mem_reg[60][35]  ( .D(n24793), .E(n6453), .CP(clk), .QN(n18031) );
  EDFD1 \Mem_reg[59][35]  ( .D(n24793), .E(n6452), .CP(clk), .QN(n4967) );
  EDFD1 \Mem_reg[58][35]  ( .D(n24793), .E(n6451), .CP(clk), .QN(n4919) );
  EDFD1 \Mem_reg[57][35]  ( .D(n24793), .E(n6450), .CP(clk), .QN(n4871) );
  EDFD1 \Mem_reg[56][35]  ( .D(n24793), .E(n6449), .CP(clk), .QN(n4823) );
  EDFD1 \Mem_reg[55][35]  ( .D(n24793), .E(n6448), .CP(clk), .QN(n4775) );
  EDFD1 \Mem_reg[54][35]  ( .D(n24793), .E(n6447), .CP(clk), .QN(n15588) );
  EDFD1 \Mem_reg[53][35]  ( .D(n24793), .E(n6446), .CP(clk), .QN(n4679) );
  EDFD1 \Mem_reg[52][35]  ( .D(n24793), .E(n6445), .CP(clk), .Q(n27176) );
  EDFD1 \Mem_reg[51][35]  ( .D(n24793), .E(n6444), .CP(clk), .QN(n4583) );
  EDFD1 \Mem_reg[50][35]  ( .D(n24793), .E(n6443), .CP(clk), .QN(n4535) );
  EDFD1 \Mem_reg[49][35]  ( .D(n24793), .E(n6442), .CP(clk), .QN(n4487) );
  EDFD1 \Mem_reg[48][35]  ( .D(n24793), .E(n6441), .CP(clk), .QN(n4439) );
  EDFD1 \Mem_reg[47][35]  ( .D(n24793), .E(n6440), .CP(clk), .QN(n4391) );
  EDFD1 \Mem_reg[46][35]  ( .D(n24793), .E(n6439), .CP(clk), .QN(n4343) );
  EDFD1 \Mem_reg[43][35]  ( .D(n24793), .E(n6438), .CP(clk), .QN(n4295) );
  EDFD1 \Mem_reg[42][35]  ( .D(n24793), .E(n6437), .CP(clk), .QN(n4247) );
  EDFD1 \Mem_reg[41][35]  ( .D(n24793), .E(n6436), .CP(clk), .QN(n4199) );
  EDFD1 \Mem_reg[40][35]  ( .D(n24793), .E(n6435), .CP(clk), .QN(n4151) );
  EDFD1 \Mem_reg[39][35]  ( .D(n24793), .E(n6434), .CP(clk), .QN(n4103) );
  EDFD1 \Mem_reg[38][35]  ( .D(n24793), .E(n6433), .CP(clk), .QN(n4055) );
  EDFD1 \Mem_reg[37][35]  ( .D(n24793), .E(n6432), .CP(clk), .QN(n4007) );
  EDFD1 \Mem_reg[36][35]  ( .D(n24793), .E(n6431), .CP(clk), .QN(n3959) );
  EDFD1 \Mem_reg[35][35]  ( .D(n24793), .E(n6430), .CP(clk), .QN(n3911) );
  EDFD1 \Mem_reg[34][35]  ( .D(n24793), .E(n6429), .CP(clk), .QN(n3863) );
  EDFD1 \Mem_reg[33][35]  ( .D(n24793), .E(n6428), .CP(clk), .QN(n3815) );
  EDFD1 \Mem_reg[32][35]  ( .D(n24793), .E(n6427), .CP(clk), .QN(n3767) );
  EDFD1 \Mem_reg[31][35]  ( .D(n24793), .E(n6426), .CP(clk), .QN(n3719) );
  EDFD1 \Mem_reg[30][35]  ( .D(n24793), .E(n6425), .CP(clk), .QN(n3671) );
  EDFD1 \Mem_reg[29][35]  ( .D(n24793), .E(n6424), .CP(clk), .QN(n3623) );
  EDFD1 \Mem_reg[28][35]  ( .D(n24793), .E(n6423), .CP(clk), .QN(n3575) );
  EDFD1 \Mem_reg[27][35]  ( .D(n24793), .E(n6422), .CP(clk), .QN(n3527) );
  EDFD1 \Mem_reg[26][35]  ( .D(n24793), .E(n6421), .CP(clk), .QN(n3479) );
  EDFD1 \Mem_reg[25][35]  ( .D(n24793), .E(n6420), .CP(clk), .QN(n3431) );
  EDFD1 \Mem_reg[24][35]  ( .D(n24793), .E(n6463), .CP(clk), .QN(n3383) );
  EDFD1 \Mem_reg[23][35]  ( .D(n24793), .E(n6464), .CP(clk), .QN(n3335) );
  EDFD1 \Mem_reg[22][35]  ( .D(n24793), .E(n6465), .CP(clk), .QN(n3287) );
  EDFD1 \Mem_reg[21][35]  ( .D(n24793), .E(n6466), .CP(clk), .QN(n3239) );
  EDFD1 \Mem_reg[20][35]  ( .D(n24793), .E(n6467), .CP(clk), .QN(n3191) );
  EDFD1 \Mem_reg[19][35]  ( .D(n24793), .E(n6468), .CP(clk), .QN(n3143) );
  EDFD1 \Mem_reg[18][35]  ( .D(n24793), .E(n6469), .CP(clk), .QN(n3095) );
  EDFD1 \Mem_reg[17][35]  ( .D(n24793), .E(n6470), .CP(clk), .QN(n3047) );
  EDFD1 \Mem_reg[16][35]  ( .D(n24793), .E(n6471), .CP(clk), .QN(n2999) );
  EDFD1 \Mem_reg[15][35]  ( .D(n24793), .E(n6472), .CP(clk), .QN(n2951) );
  EDFD1 \Mem_reg[14][35]  ( .D(n24793), .E(n24720), .CP(clk), .QN(n2903) );
  EDFD1 \Mem_reg[13][35]  ( .D(n24793), .E(n24709), .CP(clk), .QN(n2855) );
  EDFD1 \Mem_reg[12][35]  ( .D(n24793), .E(n24717), .CP(clk), .QN(n2807) );
  EDFD1 \Mem_reg[11][35]  ( .D(n24793), .E(n24707), .CP(clk), .QN(n2759) );
  EDFD1 \Mem_reg[10][35]  ( .D(n24793), .E(n6477), .CP(clk), .QN(n2711) );
  EDFD1 \Mem_reg[9][35]  ( .D(n24793), .E(n24708), .CP(clk), .QN(n2663) );
  EDFD1 \Mem_reg[8][35]  ( .D(n24793), .E(n15642), .CP(clk), .QN(n2615) );
  EDFD1 \Mem_reg[7][35]  ( .D(n24793), .E(n24718), .CP(clk), .QN(n2567) );
  EDFD1 \Mem_reg[6][35]  ( .D(n24793), .E(n24716), .CP(clk), .QN(n2519) );
  EDFD1 \Mem_reg[5][35]  ( .D(n24793), .E(n24719), .CP(clk), .QN(n2471) );
  EDFD1 \Mem_reg[4][35]  ( .D(n24793), .E(n24706), .CP(clk), .QN(n2423) );
  EDFD1 \Mem_reg[3][35]  ( .D(n24793), .E(n24721), .CP(clk), .QN(n2375) );
  EDFD1 \Mem_reg[2][35]  ( .D(n24793), .E(n6460), .CP(clk), .QN(n2327) );
  EDFD1 \Mem_reg[1][35]  ( .D(n24793), .E(n24703), .CP(clk), .QN(n2279) );
  EDFD1 \Mem_reg[0][35]  ( .D(n24793), .E(n24705), .CP(clk), .QN(n2231) );
  EDFD1 \Mem_reg[88][34]  ( .D(n24791), .E(n6419), .CP(clk), .Q(n27173) );
  EDFD1 \Mem_reg[87][34]  ( .D(n24791), .E(n6418), .CP(clk), .QN(n6312) );
  EDFD1 \Mem_reg[86][34]  ( .D(n24791), .E(n6417), .CP(clk), .QN(n24661) );
  EDFD1 \Mem_reg[85][34]  ( .D(n24791), .E(n6416), .CP(clk), .QN(n6216) );
  EDFD1 \Mem_reg[84][34]  ( .D(n24791), .E(n6415), .CP(clk), .QN(n6168) );
  EDFD1 \Mem_reg[83][34]  ( .D(n24791), .E(n6414), .CP(clk), .QN(n6120) );
  EDFD1 \Mem_reg[82][34]  ( .D(n24791), .E(n6413), .CP(clk), .QN(n6072) );
  EDFD1 \Mem_reg[81][34]  ( .D(n24791), .E(n6412), .CP(clk), .QN(n6024) );
  EDFD1 \Mem_reg[80][34]  ( .D(n24791), .E(n6411), .CP(clk), .QN(n5976) );
  EDFD1 \Mem_reg[79][34]  ( .D(n24791), .E(n6410), .CP(clk), .QN(n5928) );
  EDFD1 \Mem_reg[78][34]  ( .D(n24791), .E(n6409), .CP(clk), .QN(n5880) );
  EDFD1 \Mem_reg[77][34]  ( .D(n24791), .E(n6408), .CP(clk), .QN(n5832) );
  EDFD1 \Mem_reg[76][34]  ( .D(n24791), .E(n6407), .CP(clk), .QN(n5784) );
  EDFD1 \Mem_reg[75][34]  ( .D(n24791), .E(n6406), .CP(clk), .QN(n27174) );
  EDFD1 \Mem_reg[74][34]  ( .D(n24791), .E(n6405), .CP(clk), .QN(n5688) );
  EDFD1 \Mem_reg[73][34]  ( .D(n24791), .E(n6404), .CP(clk), .QN(n27175) );
  EDFD1 \Mem_reg[72][34]  ( .D(n24791), .E(n6403), .CP(clk), .QN(n5592) );
  EDFD1 \Mem_reg[71][34]  ( .D(n24791), .E(n6402), .CP(clk), .QN(n5544) );
  EDFD1 \Mem_reg[70][34]  ( .D(n24791), .E(n6401), .CP(clk), .QN(n5496) );
  EDFD1 \Mem_reg[69][34]  ( .D(n24791), .E(n6400), .CP(clk), .QN(n5448) );
  EDFD1 \Mem_reg[68][34]  ( .D(n24791), .E(n6399), .CP(clk), .QN(n5400) );
  EDFD1 \Mem_reg[67][34]  ( .D(n24791), .E(n6398), .CP(clk), .QN(n5352) );
  EDFD1 \Mem_reg[66][34]  ( .D(n24791), .E(n6397), .CP(clk), .QN(n5304) );
  EDFD1 \Mem_reg[65][34]  ( .D(n24791), .E(n6396), .CP(clk), .QN(n15585) );
  EDFD1 \Mem_reg[64][34]  ( .D(n24791), .E(n6395), .CP(clk), .QN(n5208) );
  EDFD1 \Mem_reg[63][34]  ( .D(n24791), .E(n6456), .CP(clk), .QN(n5160) );
  EDFD1 \Mem_reg[62][34]  ( .D(n24791), .E(n6455), .CP(clk), .QN(n5112) );
  EDFD1 \Mem_reg[61][34]  ( .D(n24791), .E(n6454), .CP(clk), .QN(n18029) );
  EDFD1 \Mem_reg[60][34]  ( .D(n24791), .E(n6453), .CP(clk), .QN(n18028) );
  EDFD1 \Mem_reg[59][34]  ( .D(n24791), .E(n6452), .CP(clk), .QN(n4968) );
  EDFD1 \Mem_reg[58][34]  ( .D(n24791), .E(n6451), .CP(clk), .QN(n4920) );
  EDFD1 \Mem_reg[57][34]  ( .D(n24791), .E(n6450), .CP(clk), .QN(n4872) );
  EDFD1 \Mem_reg[56][34]  ( .D(n24791), .E(n6449), .CP(clk), .QN(n4824) );
  EDFD1 \Mem_reg[55][34]  ( .D(n24791), .E(n6448), .CP(clk), .QN(n4776) );
  EDFD1 \Mem_reg[54][34]  ( .D(n24791), .E(n6447), .CP(clk), .QN(n15584) );
  EDFD1 \Mem_reg[53][34]  ( .D(n24791), .E(n6446), .CP(clk), .QN(n4680) );
  EDFD1 \Mem_reg[52][34]  ( .D(n24791), .E(n6445), .CP(clk), .Q(n27172) );
  EDFD1 \Mem_reg[51][34]  ( .D(n24791), .E(n6444), .CP(clk), .QN(n4584) );
  EDFD1 \Mem_reg[50][34]  ( .D(n24791), .E(n6443), .CP(clk), .QN(n4536) );
  EDFD1 \Mem_reg[49][34]  ( .D(n24791), .E(n6442), .CP(clk), .QN(n4488) );
  EDFD1 \Mem_reg[48][34]  ( .D(n24791), .E(n6441), .CP(clk), .QN(n4440) );
  EDFD1 \Mem_reg[47][34]  ( .D(n24791), .E(n6440), .CP(clk), .QN(n4392) );
  EDFD1 \Mem_reg[46][34]  ( .D(n24791), .E(n6439), .CP(clk), .QN(n4344) );
  EDFD1 \Mem_reg[43][34]  ( .D(n24791), .E(n6438), .CP(clk), .QN(n4296) );
  EDFD1 \Mem_reg[42][34]  ( .D(n24791), .E(n6437), .CP(clk), .QN(n4248) );
  EDFD1 \Mem_reg[41][34]  ( .D(n24791), .E(n6436), .CP(clk), .QN(n4200) );
  EDFD1 \Mem_reg[40][34]  ( .D(n24791), .E(n6435), .CP(clk), .QN(n4152) );
  EDFD1 \Mem_reg[39][34]  ( .D(n24791), .E(n6434), .CP(clk), .QN(n4104) );
  EDFD1 \Mem_reg[38][34]  ( .D(n24791), .E(n6433), .CP(clk), .QN(n4056) );
  EDFD1 \Mem_reg[37][34]  ( .D(n24791), .E(n6432), .CP(clk), .QN(n4008) );
  EDFD1 \Mem_reg[36][34]  ( .D(n24791), .E(n6431), .CP(clk), .QN(n3960) );
  EDFD1 \Mem_reg[35][34]  ( .D(n24791), .E(n6430), .CP(clk), .QN(n3912) );
  EDFD1 \Mem_reg[34][34]  ( .D(n24791), .E(n6429), .CP(clk), .QN(n3864) );
  EDFD1 \Mem_reg[33][34]  ( .D(n24791), .E(n6428), .CP(clk), .QN(n3816) );
  EDFD1 \Mem_reg[32][34]  ( .D(n24791), .E(n6427), .CP(clk), .QN(n3768) );
  EDFD1 \Mem_reg[31][34]  ( .D(n24791), .E(n6426), .CP(clk), .QN(n3720) );
  EDFD1 \Mem_reg[30][34]  ( .D(n24791), .E(n6425), .CP(clk), .QN(n3672) );
  EDFD1 \Mem_reg[29][34]  ( .D(n24791), .E(n6424), .CP(clk), .QN(n3624) );
  EDFD1 \Mem_reg[28][34]  ( .D(n24791), .E(n6423), .CP(clk), .QN(n3576) );
  EDFD1 \Mem_reg[27][34]  ( .D(n24791), .E(n6422), .CP(clk), .QN(n3528) );
  EDFD1 \Mem_reg[26][34]  ( .D(n24791), .E(n6421), .CP(clk), .QN(n3480) );
  EDFD1 \Mem_reg[25][34]  ( .D(n24791), .E(n6420), .CP(clk), .QN(n3432) );
  EDFD1 \Mem_reg[24][34]  ( .D(n24791), .E(n6463), .CP(clk), .QN(n3384) );
  EDFD1 \Mem_reg[23][34]  ( .D(n24791), .E(n6464), .CP(clk), .QN(n3336) );
  EDFD1 \Mem_reg[22][34]  ( .D(n24791), .E(n6465), .CP(clk), .QN(n3288) );
  EDFD1 \Mem_reg[21][34]  ( .D(n24791), .E(n6466), .CP(clk), .QN(n3240) );
  EDFD1 \Mem_reg[20][34]  ( .D(n24791), .E(n6467), .CP(clk), .QN(n3192) );
  EDFD1 \Mem_reg[19][34]  ( .D(n24791), .E(n6468), .CP(clk), .QN(n3144) );
  EDFD1 \Mem_reg[18][34]  ( .D(n24791), .E(n6469), .CP(clk), .QN(n3096) );
  EDFD1 \Mem_reg[17][34]  ( .D(n24791), .E(n6470), .CP(clk), .QN(n3048) );
  EDFD1 \Mem_reg[16][34]  ( .D(n24791), .E(n6471), .CP(clk), .QN(n3000) );
  EDFD1 \Mem_reg[15][34]  ( .D(n24791), .E(n6472), .CP(clk), .QN(n2952) );
  EDFD1 \Mem_reg[14][34]  ( .D(n24791), .E(n24720), .CP(clk), .QN(n2904) );
  EDFD1 \Mem_reg[13][34]  ( .D(n24791), .E(n24709), .CP(clk), .QN(n2856) );
  EDFD1 \Mem_reg[12][34]  ( .D(n24791), .E(n24717), .CP(clk), .QN(n2808) );
  EDFD1 \Mem_reg[11][34]  ( .D(n24791), .E(n24707), .CP(clk), .QN(n2760) );
  EDFD1 \Mem_reg[10][34]  ( .D(n24791), .E(n6477), .CP(clk), .QN(n2712) );
  EDFD1 \Mem_reg[9][34]  ( .D(n24791), .E(n24708), .CP(clk), .QN(n2664) );
  EDFD1 \Mem_reg[8][34]  ( .D(n24791), .E(n15642), .CP(clk), .QN(n2616) );
  EDFD1 \Mem_reg[7][34]  ( .D(n24791), .E(n24718), .CP(clk), .QN(n2568) );
  EDFD1 \Mem_reg[6][34]  ( .D(n24791), .E(n24716), .CP(clk), .QN(n2520) );
  EDFD1 \Mem_reg[5][34]  ( .D(n24791), .E(n24719), .CP(clk), .QN(n2472) );
  EDFD1 \Mem_reg[4][34]  ( .D(n24791), .E(n24706), .CP(clk), .QN(n2424) );
  EDFD1 \Mem_reg[3][34]  ( .D(n24791), .E(n24721), .CP(clk), .QN(n2376) );
  EDFD1 \Mem_reg[2][34]  ( .D(n24791), .E(n6460), .CP(clk), .QN(n2328) );
  EDFD1 \Mem_reg[1][34]  ( .D(n24791), .E(n24703), .CP(clk), .QN(n2280) );
  EDFD1 \Mem_reg[0][34]  ( .D(n24791), .E(n24705), .CP(clk), .QN(n2232) );
  EDFD1 \Mem_reg[88][33]  ( .D(n24789), .E(n6419), .CP(clk), .Q(n27169) );
  EDFD1 \Mem_reg[87][33]  ( .D(n24789), .E(n6418), .CP(clk), .QN(n6313) );
  EDFD1 \Mem_reg[86][33]  ( .D(n24789), .E(n6417), .CP(clk), .QN(n24658) );
  EDFD1 \Mem_reg[85][33]  ( .D(n24789), .E(n6416), .CP(clk), .QN(n6217) );
  EDFD1 \Mem_reg[84][33]  ( .D(n24789), .E(n6415), .CP(clk), .QN(n6169) );
  EDFD1 \Mem_reg[83][33]  ( .D(n24789), .E(n6414), .CP(clk), .QN(n6121) );
  EDFD1 \Mem_reg[82][33]  ( .D(n24789), .E(n6413), .CP(clk), .QN(n6073) );
  EDFD1 \Mem_reg[81][33]  ( .D(n24789), .E(n6412), .CP(clk), .QN(n6025) );
  EDFD1 \Mem_reg[80][33]  ( .D(n24789), .E(n6411), .CP(clk), .QN(n5977) );
  EDFD1 \Mem_reg[79][33]  ( .D(n24789), .E(n6410), .CP(clk), .QN(n5929) );
  EDFD1 \Mem_reg[78][33]  ( .D(n24789), .E(n6409), .CP(clk), .QN(n5881) );
  EDFD1 \Mem_reg[77][33]  ( .D(n24789), .E(n6408), .CP(clk), .QN(n5833) );
  EDFD1 \Mem_reg[76][33]  ( .D(n24789), .E(n6407), .CP(clk), .QN(n5785) );
  EDFD1 \Mem_reg[75][33]  ( .D(n24789), .E(n6406), .CP(clk), .QN(n27170) );
  EDFD1 \Mem_reg[74][33]  ( .D(n24789), .E(n6405), .CP(clk), .QN(n5689) );
  EDFD1 \Mem_reg[73][33]  ( .D(n24789), .E(n6404), .CP(clk), .QN(n27171) );
  EDFD1 \Mem_reg[72][33]  ( .D(n24789), .E(n6403), .CP(clk), .QN(n5593) );
  EDFD1 \Mem_reg[71][33]  ( .D(n24789), .E(n6402), .CP(clk), .QN(n5545) );
  EDFD1 \Mem_reg[70][33]  ( .D(n24789), .E(n6401), .CP(clk), .QN(n5497) );
  EDFD1 \Mem_reg[69][33]  ( .D(n24789), .E(n6400), .CP(clk), .QN(n5449) );
  EDFD1 \Mem_reg[68][33]  ( .D(n24789), .E(n6399), .CP(clk), .QN(n5401) );
  EDFD1 \Mem_reg[67][33]  ( .D(n24789), .E(n6398), .CP(clk), .QN(n5353) );
  EDFD1 \Mem_reg[66][33]  ( .D(n24789), .E(n6397), .CP(clk), .QN(n5305) );
  EDFD1 \Mem_reg[65][33]  ( .D(n24789), .E(n6396), .CP(clk), .QN(n15581) );
  EDFD1 \Mem_reg[64][33]  ( .D(n24789), .E(n6395), .CP(clk), .QN(n5209) );
  EDFD1 \Mem_reg[63][33]  ( .D(n24789), .E(n6456), .CP(clk), .QN(n5161) );
  EDFD1 \Mem_reg[62][33]  ( .D(n24789), .E(n6455), .CP(clk), .QN(n5113) );
  EDFD1 \Mem_reg[61][33]  ( .D(n24789), .E(n6454), .CP(clk), .QN(n18026) );
  EDFD1 \Mem_reg[60][33]  ( .D(n24789), .E(n6453), .CP(clk), .QN(n18025) );
  EDFD1 \Mem_reg[59][33]  ( .D(n24789), .E(n6452), .CP(clk), .QN(n4969) );
  EDFD1 \Mem_reg[58][33]  ( .D(n24789), .E(n6451), .CP(clk), .QN(n4921) );
  EDFD1 \Mem_reg[57][33]  ( .D(n24789), .E(n6450), .CP(clk), .QN(n4873) );
  EDFD1 \Mem_reg[56][33]  ( .D(n24789), .E(n6449), .CP(clk), .QN(n4825) );
  EDFD1 \Mem_reg[55][33]  ( .D(n24789), .E(n6448), .CP(clk), .QN(n4777) );
  EDFD1 \Mem_reg[54][33]  ( .D(n24789), .E(n6447), .CP(clk), .QN(n15580) );
  EDFD1 \Mem_reg[53][33]  ( .D(n24789), .E(n6446), .CP(clk), .QN(n4681) );
  EDFD1 \Mem_reg[52][33]  ( .D(n24789), .E(n6445), .CP(clk), .Q(n27168) );
  EDFD1 \Mem_reg[51][33]  ( .D(n24789), .E(n6444), .CP(clk), .QN(n4585) );
  EDFD1 \Mem_reg[50][33]  ( .D(n24789), .E(n6443), .CP(clk), .QN(n4537) );
  EDFD1 \Mem_reg[49][33]  ( .D(n24789), .E(n6442), .CP(clk), .QN(n4489) );
  EDFD1 \Mem_reg[48][33]  ( .D(n24789), .E(n6441), .CP(clk), .QN(n4441) );
  EDFD1 \Mem_reg[47][33]  ( .D(n24789), .E(n6440), .CP(clk), .QN(n4393) );
  EDFD1 \Mem_reg[46][33]  ( .D(n24789), .E(n6439), .CP(clk), .QN(n4345) );
  EDFD1 \Mem_reg[43][33]  ( .D(n24789), .E(n6438), .CP(clk), .QN(n4297) );
  EDFD1 \Mem_reg[42][33]  ( .D(n24789), .E(n6437), .CP(clk), .QN(n4249) );
  EDFD1 \Mem_reg[41][33]  ( .D(n24789), .E(n6436), .CP(clk), .QN(n4201) );
  EDFD1 \Mem_reg[40][33]  ( .D(n24789), .E(n6435), .CP(clk), .QN(n4153) );
  EDFD1 \Mem_reg[39][33]  ( .D(n24789), .E(n6434), .CP(clk), .QN(n4105) );
  EDFD1 \Mem_reg[38][33]  ( .D(n24789), .E(n6433), .CP(clk), .QN(n4057) );
  EDFD1 \Mem_reg[37][33]  ( .D(n24789), .E(n6432), .CP(clk), .QN(n4009) );
  EDFD1 \Mem_reg[36][33]  ( .D(n24789), .E(n6431), .CP(clk), .QN(n3961) );
  EDFD1 \Mem_reg[35][33]  ( .D(n24789), .E(n6430), .CP(clk), .QN(n3913) );
  EDFD1 \Mem_reg[34][33]  ( .D(n24789), .E(n6429), .CP(clk), .QN(n3865) );
  EDFD1 \Mem_reg[33][33]  ( .D(n24789), .E(n6428), .CP(clk), .QN(n3817) );
  EDFD1 \Mem_reg[32][33]  ( .D(n24789), .E(n6427), .CP(clk), .QN(n3769) );
  EDFD1 \Mem_reg[31][33]  ( .D(n24789), .E(n6426), .CP(clk), .QN(n3721) );
  EDFD1 \Mem_reg[30][33]  ( .D(n24789), .E(n6425), .CP(clk), .QN(n3673) );
  EDFD1 \Mem_reg[29][33]  ( .D(n24789), .E(n6424), .CP(clk), .QN(n3625) );
  EDFD1 \Mem_reg[28][33]  ( .D(n24789), .E(n6423), .CP(clk), .QN(n3577) );
  EDFD1 \Mem_reg[27][33]  ( .D(n24789), .E(n6422), .CP(clk), .QN(n3529) );
  EDFD1 \Mem_reg[26][33]  ( .D(n24789), .E(n6421), .CP(clk), .QN(n3481) );
  EDFD1 \Mem_reg[25][33]  ( .D(n24789), .E(n6420), .CP(clk), .QN(n3433) );
  EDFD1 \Mem_reg[24][33]  ( .D(n24789), .E(n6463), .CP(clk), .QN(n3385) );
  EDFD1 \Mem_reg[23][33]  ( .D(n24789), .E(n6464), .CP(clk), .QN(n3337) );
  EDFD1 \Mem_reg[22][33]  ( .D(n24789), .E(n6465), .CP(clk), .QN(n3289) );
  EDFD1 \Mem_reg[21][33]  ( .D(n24789), .E(n6466), .CP(clk), .QN(n3241) );
  EDFD1 \Mem_reg[20][33]  ( .D(n24789), .E(n6467), .CP(clk), .QN(n3193) );
  EDFD1 \Mem_reg[19][33]  ( .D(n24789), .E(n6468), .CP(clk), .QN(n3145) );
  EDFD1 \Mem_reg[18][33]  ( .D(n24789), .E(n6469), .CP(clk), .QN(n3097) );
  EDFD1 \Mem_reg[17][33]  ( .D(n24789), .E(n6470), .CP(clk), .QN(n3049) );
  EDFD1 \Mem_reg[16][33]  ( .D(n24789), .E(n6471), .CP(clk), .QN(n3001) );
  EDFD1 \Mem_reg[15][33]  ( .D(n24789), .E(n6472), .CP(clk), .QN(n2953) );
  EDFD1 \Mem_reg[14][33]  ( .D(n24789), .E(n24720), .CP(clk), .QN(n2905) );
  EDFD1 \Mem_reg[13][33]  ( .D(n24789), .E(n24709), .CP(clk), .QN(n2857) );
  EDFD1 \Mem_reg[12][33]  ( .D(n24789), .E(n24717), .CP(clk), .QN(n2809) );
  EDFD1 \Mem_reg[11][33]  ( .D(n24789), .E(n24707), .CP(clk), .QN(n2761) );
  EDFD1 \Mem_reg[10][33]  ( .D(n24789), .E(n6477), .CP(clk), .QN(n2713) );
  EDFD1 \Mem_reg[9][33]  ( .D(n24789), .E(n24708), .CP(clk), .QN(n2665) );
  EDFD1 \Mem_reg[8][33]  ( .D(n24789), .E(n15642), .CP(clk), .QN(n2617) );
  EDFD1 \Mem_reg[7][33]  ( .D(n24789), .E(n24718), .CP(clk), .QN(n2569) );
  EDFD1 \Mem_reg[6][33]  ( .D(n24789), .E(n24716), .CP(clk), .QN(n2521) );
  EDFD1 \Mem_reg[5][33]  ( .D(n24789), .E(n24719), .CP(clk), .QN(n2473) );
  EDFD1 \Mem_reg[4][33]  ( .D(n24789), .E(n24706), .CP(clk), .QN(n2425) );
  EDFD1 \Mem_reg[3][33]  ( .D(n24789), .E(n24721), .CP(clk), .QN(n2377) );
  EDFD1 \Mem_reg[2][33]  ( .D(n24789), .E(n6460), .CP(clk), .QN(n2329) );
  EDFD1 \Mem_reg[1][33]  ( .D(n24789), .E(n24703), .CP(clk), .QN(n2281) );
  EDFD1 \Mem_reg[0][33]  ( .D(n24789), .E(n24705), .CP(clk), .QN(n2233) );
  EDFD1 \Mem_reg[88][32]  ( .D(n24787), .E(n6419), .CP(clk), .Q(n27165) );
  EDFD1 \Mem_reg[87][32]  ( .D(n24787), .E(n6418), .CP(clk), .QN(n6314) );
  EDFD1 \Mem_reg[86][32]  ( .D(n24787), .E(n6417), .CP(clk), .QN(n24655) );
  EDFD1 \Mem_reg[85][32]  ( .D(n24787), .E(n6416), .CP(clk), .QN(n6218) );
  EDFD1 \Mem_reg[84][32]  ( .D(n24787), .E(n6415), .CP(clk), .QN(n6170) );
  EDFD1 \Mem_reg[83][32]  ( .D(n24787), .E(n6414), .CP(clk), .QN(n6122) );
  EDFD1 \Mem_reg[82][32]  ( .D(n24787), .E(n6413), .CP(clk), .QN(n6074) );
  EDFD1 \Mem_reg[81][32]  ( .D(n24787), .E(n6412), .CP(clk), .QN(n6026) );
  EDFD1 \Mem_reg[80][32]  ( .D(n24787), .E(n6411), .CP(clk), .QN(n5978) );
  EDFD1 \Mem_reg[79][32]  ( .D(n24787), .E(n6410), .CP(clk), .QN(n5930) );
  EDFD1 \Mem_reg[78][32]  ( .D(n24787), .E(n6409), .CP(clk), .QN(n5882) );
  EDFD1 \Mem_reg[77][32]  ( .D(n24787), .E(n6408), .CP(clk), .QN(n5834) );
  EDFD1 \Mem_reg[76][32]  ( .D(n24787), .E(n6407), .CP(clk), .QN(n5786) );
  EDFD1 \Mem_reg[75][32]  ( .D(n24787), .E(n6406), .CP(clk), .QN(n27166) );
  EDFD1 \Mem_reg[74][32]  ( .D(n24787), .E(n6405), .CP(clk), .QN(n5690) );
  EDFD1 \Mem_reg[73][32]  ( .D(n24787), .E(n6404), .CP(clk), .QN(n27167) );
  EDFD1 \Mem_reg[72][32]  ( .D(n24787), .E(n6403), .CP(clk), .QN(n5594) );
  EDFD1 \Mem_reg[71][32]  ( .D(n24787), .E(n6402), .CP(clk), .QN(n5546) );
  EDFD1 \Mem_reg[70][32]  ( .D(n24787), .E(n6401), .CP(clk), .QN(n5498) );
  EDFD1 \Mem_reg[69][32]  ( .D(n24787), .E(n6400), .CP(clk), .QN(n5450) );
  EDFD1 \Mem_reg[68][32]  ( .D(n24787), .E(n6399), .CP(clk), .QN(n5402) );
  EDFD1 \Mem_reg[67][32]  ( .D(n24787), .E(n6398), .CP(clk), .QN(n5354) );
  EDFD1 \Mem_reg[66][32]  ( .D(n24787), .E(n6397), .CP(clk), .QN(n5306) );
  EDFD1 \Mem_reg[65][32]  ( .D(n24787), .E(n6396), .CP(clk), .QN(n15577) );
  EDFD1 \Mem_reg[64][32]  ( .D(n24787), .E(n6395), .CP(clk), .QN(n5210) );
  EDFD1 \Mem_reg[63][32]  ( .D(n24787), .E(n6456), .CP(clk), .QN(n5162) );
  EDFD1 \Mem_reg[62][32]  ( .D(n24787), .E(n6455), .CP(clk), .QN(n5114) );
  EDFD1 \Mem_reg[61][32]  ( .D(n24787), .E(n6454), .CP(clk), .QN(n18023) );
  EDFD1 \Mem_reg[60][32]  ( .D(n24787), .E(n6453), .CP(clk), .QN(n18022) );
  EDFD1 \Mem_reg[59][32]  ( .D(n24787), .E(n6452), .CP(clk), .QN(n4970) );
  EDFD1 \Mem_reg[58][32]  ( .D(n24787), .E(n6451), .CP(clk), .QN(n4922) );
  EDFD1 \Mem_reg[57][32]  ( .D(n24787), .E(n6450), .CP(clk), .QN(n4874) );
  EDFD1 \Mem_reg[56][32]  ( .D(n24787), .E(n6449), .CP(clk), .QN(n4826) );
  EDFD1 \Mem_reg[55][32]  ( .D(n24787), .E(n6448), .CP(clk), .QN(n4778) );
  EDFD1 \Mem_reg[54][32]  ( .D(n24787), .E(n6447), .CP(clk), .QN(n15576) );
  EDFD1 \Mem_reg[53][32]  ( .D(n24787), .E(n6446), .CP(clk), .QN(n4682) );
  EDFD1 \Mem_reg[52][32]  ( .D(n24787), .E(n6445), .CP(clk), .Q(n27164) );
  EDFD1 \Mem_reg[51][32]  ( .D(n24787), .E(n6444), .CP(clk), .QN(n4586) );
  EDFD1 \Mem_reg[50][32]  ( .D(n24787), .E(n6443), .CP(clk), .QN(n4538) );
  EDFD1 \Mem_reg[49][32]  ( .D(n24787), .E(n6442), .CP(clk), .QN(n4490) );
  EDFD1 \Mem_reg[48][32]  ( .D(n24787), .E(n6441), .CP(clk), .QN(n4442) );
  EDFD1 \Mem_reg[47][32]  ( .D(n24787), .E(n6440), .CP(clk), .QN(n4394) );
  EDFD1 \Mem_reg[46][32]  ( .D(n24787), .E(n6439), .CP(clk), .QN(n4346) );
  EDFD1 \Mem_reg[43][32]  ( .D(n24787), .E(n6438), .CP(clk), .QN(n4298) );
  EDFD1 \Mem_reg[42][32]  ( .D(n24787), .E(n6437), .CP(clk), .QN(n4250) );
  EDFD1 \Mem_reg[41][32]  ( .D(n24787), .E(n6436), .CP(clk), .QN(n4202) );
  EDFD1 \Mem_reg[40][32]  ( .D(n24787), .E(n6435), .CP(clk), .QN(n4154) );
  EDFD1 \Mem_reg[39][32]  ( .D(n24787), .E(n6434), .CP(clk), .QN(n4106) );
  EDFD1 \Mem_reg[38][32]  ( .D(n24787), .E(n6433), .CP(clk), .QN(n4058) );
  EDFD1 \Mem_reg[37][32]  ( .D(n24787), .E(n6432), .CP(clk), .QN(n4010) );
  EDFD1 \Mem_reg[36][32]  ( .D(n24787), .E(n6431), .CP(clk), .QN(n3962) );
  EDFD1 \Mem_reg[35][32]  ( .D(n24787), .E(n6430), .CP(clk), .QN(n3914) );
  EDFD1 \Mem_reg[34][32]  ( .D(n24787), .E(n6429), .CP(clk), .QN(n3866) );
  EDFD1 \Mem_reg[33][32]  ( .D(n24787), .E(n6428), .CP(clk), .QN(n3818) );
  EDFD1 \Mem_reg[32][32]  ( .D(n24787), .E(n6427), .CP(clk), .QN(n3770) );
  EDFD1 \Mem_reg[31][32]  ( .D(n24787), .E(n6426), .CP(clk), .QN(n3722) );
  EDFD1 \Mem_reg[30][32]  ( .D(n24787), .E(n6425), .CP(clk), .QN(n3674) );
  EDFD1 \Mem_reg[29][32]  ( .D(n24787), .E(n6424), .CP(clk), .QN(n3626) );
  EDFD1 \Mem_reg[28][32]  ( .D(n24787), .E(n6423), .CP(clk), .QN(n3578) );
  EDFD1 \Mem_reg[27][32]  ( .D(n24787), .E(n6422), .CP(clk), .QN(n3530) );
  EDFD1 \Mem_reg[26][32]  ( .D(n24787), .E(n6421), .CP(clk), .QN(n3482) );
  EDFD1 \Mem_reg[25][32]  ( .D(n24787), .E(n6420), .CP(clk), .QN(n3434) );
  EDFD1 \Mem_reg[24][32]  ( .D(n24787), .E(n6463), .CP(clk), .QN(n3386) );
  EDFD1 \Mem_reg[23][32]  ( .D(n24787), .E(n6464), .CP(clk), .QN(n3338) );
  EDFD1 \Mem_reg[22][32]  ( .D(n24787), .E(n6465), .CP(clk), .QN(n3290) );
  EDFD1 \Mem_reg[21][32]  ( .D(n24787), .E(n6466), .CP(clk), .QN(n3242) );
  EDFD1 \Mem_reg[20][32]  ( .D(n24787), .E(n6467), .CP(clk), .QN(n3194) );
  EDFD1 \Mem_reg[19][32]  ( .D(n24787), .E(n6468), .CP(clk), .QN(n3146) );
  EDFD1 \Mem_reg[18][32]  ( .D(n24787), .E(n6469), .CP(clk), .QN(n3098) );
  EDFD1 \Mem_reg[17][32]  ( .D(n24787), .E(n6470), .CP(clk), .QN(n3050) );
  EDFD1 \Mem_reg[16][32]  ( .D(n24787), .E(n6471), .CP(clk), .QN(n3002) );
  EDFD1 \Mem_reg[15][32]  ( .D(n24787), .E(n6472), .CP(clk), .QN(n2954) );
  EDFD1 \Mem_reg[14][32]  ( .D(n24787), .E(n24720), .CP(clk), .QN(n2906) );
  EDFD1 \Mem_reg[13][32]  ( .D(n24787), .E(n24709), .CP(clk), .QN(n2858) );
  EDFD1 \Mem_reg[12][32]  ( .D(n24787), .E(n24717), .CP(clk), .QN(n2810) );
  EDFD1 \Mem_reg[11][32]  ( .D(n24787), .E(n24707), .CP(clk), .QN(n2762) );
  EDFD1 \Mem_reg[10][32]  ( .D(n24787), .E(n6477), .CP(clk), .QN(n2714) );
  EDFD1 \Mem_reg[9][32]  ( .D(n24787), .E(n24708), .CP(clk), .QN(n2666) );
  EDFD1 \Mem_reg[8][32]  ( .D(n24787), .E(n15642), .CP(clk), .QN(n2618) );
  EDFD1 \Mem_reg[7][32]  ( .D(n24787), .E(n24718), .CP(clk), .QN(n2570) );
  EDFD1 \Mem_reg[6][32]  ( .D(n24787), .E(n24716), .CP(clk), .QN(n2522) );
  EDFD1 \Mem_reg[5][32]  ( .D(n24787), .E(n24719), .CP(clk), .QN(n2474) );
  EDFD1 \Mem_reg[4][32]  ( .D(n24787), .E(n24706), .CP(clk), .QN(n2426) );
  EDFD1 \Mem_reg[3][32]  ( .D(n24787), .E(n24721), .CP(clk), .QN(n2378) );
  EDFD1 \Mem_reg[2][32]  ( .D(n24787), .E(n6460), .CP(clk), .QN(n2330) );
  EDFD1 \Mem_reg[1][32]  ( .D(n24787), .E(n24703), .CP(clk), .QN(n2282) );
  EDFD1 \Mem_reg[0][32]  ( .D(n24787), .E(n24705), .CP(clk), .QN(n2234) );
  EDFD1 \Mem_reg[88][31]  ( .D(n24785), .E(n6419), .CP(clk), .Q(n27161) );
  EDFD1 \Mem_reg[87][31]  ( .D(n24785), .E(n6418), .CP(clk), .QN(n6315) );
  EDFD1 \Mem_reg[86][31]  ( .D(n24785), .E(n6417), .CP(clk), .QN(n24652) );
  EDFD1 \Mem_reg[85][31]  ( .D(n24785), .E(n6416), .CP(clk), .QN(n6219) );
  EDFD1 \Mem_reg[84][31]  ( .D(n24785), .E(n6415), .CP(clk), .QN(n6171) );
  EDFD1 \Mem_reg[83][31]  ( .D(n24785), .E(n6414), .CP(clk), .QN(n6123) );
  EDFD1 \Mem_reg[82][31]  ( .D(n24785), .E(n6413), .CP(clk), .QN(n6075) );
  EDFD1 \Mem_reg[81][31]  ( .D(n24785), .E(n6412), .CP(clk), .QN(n6027) );
  EDFD1 \Mem_reg[80][31]  ( .D(n24785), .E(n6411), .CP(clk), .QN(n5979) );
  EDFD1 \Mem_reg[79][31]  ( .D(n24785), .E(n6410), .CP(clk), .QN(n5931) );
  EDFD1 \Mem_reg[78][31]  ( .D(n24785), .E(n6409), .CP(clk), .QN(n5883) );
  EDFD1 \Mem_reg[77][31]  ( .D(n24785), .E(n6408), .CP(clk), .QN(n5835) );
  EDFD1 \Mem_reg[76][31]  ( .D(n24785), .E(n6407), .CP(clk), .QN(n5787) );
  EDFD1 \Mem_reg[75][31]  ( .D(n24785), .E(n6406), .CP(clk), .QN(n27162) );
  EDFD1 \Mem_reg[74][31]  ( .D(n24785), .E(n6405), .CP(clk), .QN(n5691) );
  EDFD1 \Mem_reg[73][31]  ( .D(n24785), .E(n6404), .CP(clk), .QN(n27163) );
  EDFD1 \Mem_reg[72][31]  ( .D(n24785), .E(n6403), .CP(clk), .QN(n5595) );
  EDFD1 \Mem_reg[71][31]  ( .D(n24785), .E(n6402), .CP(clk), .QN(n5547) );
  EDFD1 \Mem_reg[70][31]  ( .D(n24785), .E(n6401), .CP(clk), .QN(n5499) );
  EDFD1 \Mem_reg[69][31]  ( .D(n24785), .E(n6400), .CP(clk), .QN(n5451) );
  EDFD1 \Mem_reg[68][31]  ( .D(n24785), .E(n6399), .CP(clk), .QN(n5403) );
  EDFD1 \Mem_reg[67][31]  ( .D(n24785), .E(n6398), .CP(clk), .QN(n5355) );
  EDFD1 \Mem_reg[66][31]  ( .D(n24785), .E(n6397), .CP(clk), .QN(n5307) );
  EDFD1 \Mem_reg[65][31]  ( .D(n24785), .E(n6396), .CP(clk), .QN(n15573) );
  EDFD1 \Mem_reg[64][31]  ( .D(n24785), .E(n6395), .CP(clk), .QN(n5211) );
  EDFD1 \Mem_reg[63][31]  ( .D(n24785), .E(n6456), .CP(clk), .QN(n5163) );
  EDFD1 \Mem_reg[62][31]  ( .D(n24785), .E(n6455), .CP(clk), .QN(n5115) );
  EDFD1 \Mem_reg[61][31]  ( .D(n24785), .E(n6454), .CP(clk), .QN(n18020) );
  EDFD1 \Mem_reg[60][31]  ( .D(n24785), .E(n6453), .CP(clk), .QN(n18019) );
  EDFD1 \Mem_reg[59][31]  ( .D(n24785), .E(n6452), .CP(clk), .QN(n4971) );
  EDFD1 \Mem_reg[58][31]  ( .D(n24785), .E(n6451), .CP(clk), .QN(n4923) );
  EDFD1 \Mem_reg[57][31]  ( .D(n24785), .E(n6450), .CP(clk), .QN(n4875) );
  EDFD1 \Mem_reg[56][31]  ( .D(n24785), .E(n6449), .CP(clk), .QN(n4827) );
  EDFD1 \Mem_reg[55][31]  ( .D(n24785), .E(n6448), .CP(clk), .QN(n4779) );
  EDFD1 \Mem_reg[54][31]  ( .D(n24785), .E(n6447), .CP(clk), .QN(n15572) );
  EDFD1 \Mem_reg[53][31]  ( .D(n24785), .E(n6446), .CP(clk), .QN(n4683) );
  EDFD1 \Mem_reg[52][31]  ( .D(n24785), .E(n6445), .CP(clk), .Q(n27160) );
  EDFD1 \Mem_reg[51][31]  ( .D(n24785), .E(n6444), .CP(clk), .QN(n4587) );
  EDFD1 \Mem_reg[50][31]  ( .D(n24785), .E(n6443), .CP(clk), .QN(n4539) );
  EDFD1 \Mem_reg[49][31]  ( .D(n24785), .E(n6442), .CP(clk), .QN(n4491) );
  EDFD1 \Mem_reg[48][31]  ( .D(n24785), .E(n6441), .CP(clk), .QN(n4443) );
  EDFD1 \Mem_reg[47][31]  ( .D(n24785), .E(n6440), .CP(clk), .QN(n4395) );
  EDFD1 \Mem_reg[46][31]  ( .D(n24785), .E(n6439), .CP(clk), .QN(n4347) );
  EDFD1 \Mem_reg[43][31]  ( .D(n24785), .E(n6438), .CP(clk), .QN(n4299) );
  EDFD1 \Mem_reg[42][31]  ( .D(n24785), .E(n6437), .CP(clk), .QN(n4251) );
  EDFD1 \Mem_reg[41][31]  ( .D(n24785), .E(n6436), .CP(clk), .QN(n4203) );
  EDFD1 \Mem_reg[40][31]  ( .D(n24785), .E(n6435), .CP(clk), .QN(n4155) );
  EDFD1 \Mem_reg[39][31]  ( .D(n24785), .E(n6434), .CP(clk), .QN(n4107) );
  EDFD1 \Mem_reg[38][31]  ( .D(n24785), .E(n6433), .CP(clk), .QN(n4059) );
  EDFD1 \Mem_reg[37][31]  ( .D(n24785), .E(n6432), .CP(clk), .QN(n4011) );
  EDFD1 \Mem_reg[36][31]  ( .D(n24785), .E(n6431), .CP(clk), .QN(n3963) );
  EDFD1 \Mem_reg[35][31]  ( .D(n24785), .E(n6430), .CP(clk), .QN(n3915) );
  EDFD1 \Mem_reg[34][31]  ( .D(n24785), .E(n6429), .CP(clk), .QN(n3867) );
  EDFD1 \Mem_reg[33][31]  ( .D(n24785), .E(n6428), .CP(clk), .QN(n3819) );
  EDFD1 \Mem_reg[32][31]  ( .D(n24785), .E(n6427), .CP(clk), .QN(n3771) );
  EDFD1 \Mem_reg[31][31]  ( .D(n24785), .E(n6426), .CP(clk), .QN(n3723) );
  EDFD1 \Mem_reg[30][31]  ( .D(n24785), .E(n6425), .CP(clk), .QN(n3675) );
  EDFD1 \Mem_reg[29][31]  ( .D(n24785), .E(n6424), .CP(clk), .QN(n3627) );
  EDFD1 \Mem_reg[28][31]  ( .D(n24785), .E(n6423), .CP(clk), .QN(n3579) );
  EDFD1 \Mem_reg[27][31]  ( .D(n24785), .E(n6422), .CP(clk), .QN(n3531) );
  EDFD1 \Mem_reg[26][31]  ( .D(n24785), .E(n6421), .CP(clk), .QN(n3483) );
  EDFD1 \Mem_reg[25][31]  ( .D(n24785), .E(n6420), .CP(clk), .QN(n3435) );
  EDFD1 \Mem_reg[24][31]  ( .D(n24785), .E(n6463), .CP(clk), .QN(n3387) );
  EDFD1 \Mem_reg[23][31]  ( .D(n24785), .E(n6464), .CP(clk), .QN(n3339) );
  EDFD1 \Mem_reg[22][31]  ( .D(n24785), .E(n6465), .CP(clk), .QN(n3291) );
  EDFD1 \Mem_reg[21][31]  ( .D(n24785), .E(n6466), .CP(clk), .QN(n3243) );
  EDFD1 \Mem_reg[20][31]  ( .D(n24785), .E(n6467), .CP(clk), .QN(n3195) );
  EDFD1 \Mem_reg[19][31]  ( .D(n24785), .E(n6468), .CP(clk), .QN(n3147) );
  EDFD1 \Mem_reg[18][31]  ( .D(n24785), .E(n6469), .CP(clk), .QN(n3099) );
  EDFD1 \Mem_reg[17][31]  ( .D(n24785), .E(n6470), .CP(clk), .QN(n3051) );
  EDFD1 \Mem_reg[16][31]  ( .D(n24785), .E(n6471), .CP(clk), .QN(n3003) );
  EDFD1 \Mem_reg[15][31]  ( .D(n24785), .E(n6472), .CP(clk), .QN(n2955) );
  EDFD1 \Mem_reg[14][31]  ( .D(n24785), .E(n24720), .CP(clk), .QN(n2907) );
  EDFD1 \Mem_reg[13][31]  ( .D(n24785), .E(n24709), .CP(clk), .QN(n2859) );
  EDFD1 \Mem_reg[12][31]  ( .D(n24785), .E(n24717), .CP(clk), .QN(n2811) );
  EDFD1 \Mem_reg[11][31]  ( .D(n24785), .E(n24707), .CP(clk), .QN(n2763) );
  EDFD1 \Mem_reg[10][31]  ( .D(n24785), .E(n6477), .CP(clk), .QN(n2715) );
  EDFD1 \Mem_reg[9][31]  ( .D(n24785), .E(n24708), .CP(clk), .QN(n2667) );
  EDFD1 \Mem_reg[8][31]  ( .D(n24785), .E(n15642), .CP(clk), .QN(n2619) );
  EDFD1 \Mem_reg[7][31]  ( .D(n24785), .E(n24718), .CP(clk), .QN(n2571) );
  EDFD1 \Mem_reg[6][31]  ( .D(n24785), .E(n24716), .CP(clk), .QN(n2523) );
  EDFD1 \Mem_reg[5][31]  ( .D(n24785), .E(n24719), .CP(clk), .QN(n2475) );
  EDFD1 \Mem_reg[4][31]  ( .D(n24785), .E(n24706), .CP(clk), .QN(n2427) );
  EDFD1 \Mem_reg[3][31]  ( .D(n24785), .E(n24721), .CP(clk), .QN(n2379) );
  EDFD1 \Mem_reg[2][31]  ( .D(n24785), .E(n6460), .CP(clk), .QN(n2331) );
  EDFD1 \Mem_reg[1][31]  ( .D(n24785), .E(n24703), .CP(clk), .QN(n2283) );
  EDFD1 \Mem_reg[0][31]  ( .D(n24785), .E(n24705), .CP(clk), .QN(n2235) );
  EDFD1 \Mem_reg[88][30]  ( .D(n24783), .E(n6419), .CP(clk), .Q(n27157) );
  EDFD1 \Mem_reg[87][30]  ( .D(n24783), .E(n6418), .CP(clk), .QN(n6316) );
  EDFD1 \Mem_reg[86][30]  ( .D(n24783), .E(n6417), .CP(clk), .QN(n24649) );
  EDFD1 \Mem_reg[85][30]  ( .D(n24783), .E(n6416), .CP(clk), .QN(n6220) );
  EDFD1 \Mem_reg[84][30]  ( .D(n24783), .E(n6415), .CP(clk), .QN(n6172) );
  EDFD1 \Mem_reg[83][30]  ( .D(n24783), .E(n6414), .CP(clk), .QN(n6124) );
  EDFD1 \Mem_reg[82][30]  ( .D(n24783), .E(n6413), .CP(clk), .QN(n6076) );
  EDFD1 \Mem_reg[81][30]  ( .D(n24783), .E(n6412), .CP(clk), .QN(n6028) );
  EDFD1 \Mem_reg[80][30]  ( .D(n24783), .E(n6411), .CP(clk), .QN(n5980) );
  EDFD1 \Mem_reg[79][30]  ( .D(n24783), .E(n6410), .CP(clk), .QN(n5932) );
  EDFD1 \Mem_reg[78][30]  ( .D(n24783), .E(n6409), .CP(clk), .QN(n5884) );
  EDFD1 \Mem_reg[77][30]  ( .D(n24783), .E(n6408), .CP(clk), .QN(n5836) );
  EDFD1 \Mem_reg[76][30]  ( .D(n24783), .E(n6407), .CP(clk), .QN(n5788) );
  EDFD1 \Mem_reg[75][30]  ( .D(n24783), .E(n6406), .CP(clk), .QN(n27158) );
  EDFD1 \Mem_reg[74][30]  ( .D(n24783), .E(n6405), .CP(clk), .QN(n5692) );
  EDFD1 \Mem_reg[73][30]  ( .D(n24783), .E(n6404), .CP(clk), .QN(n27159) );
  EDFD1 \Mem_reg[72][30]  ( .D(n24783), .E(n6403), .CP(clk), .QN(n5596) );
  EDFD1 \Mem_reg[71][30]  ( .D(n24783), .E(n6402), .CP(clk), .QN(n5548) );
  EDFD1 \Mem_reg[70][30]  ( .D(n24783), .E(n6401), .CP(clk), .QN(n5500) );
  EDFD1 \Mem_reg[69][30]  ( .D(n24783), .E(n6400), .CP(clk), .QN(n5452) );
  EDFD1 \Mem_reg[68][30]  ( .D(n24783), .E(n6399), .CP(clk), .QN(n5404) );
  EDFD1 \Mem_reg[67][30]  ( .D(n24783), .E(n6398), .CP(clk), .QN(n5356) );
  EDFD1 \Mem_reg[66][30]  ( .D(n24783), .E(n6397), .CP(clk), .QN(n5308) );
  EDFD1 \Mem_reg[65][30]  ( .D(n24783), .E(n6396), .CP(clk), .QN(n15569) );
  EDFD1 \Mem_reg[64][30]  ( .D(n24783), .E(n6395), .CP(clk), .QN(n5212) );
  EDFD1 \Mem_reg[63][30]  ( .D(n24783), .E(n6456), .CP(clk), .QN(n5164) );
  EDFD1 \Mem_reg[62][30]  ( .D(n24783), .E(n6455), .CP(clk), .QN(n5116) );
  EDFD1 \Mem_reg[61][30]  ( .D(n24783), .E(n6454), .CP(clk), .QN(n18017) );
  EDFD1 \Mem_reg[60][30]  ( .D(n24783), .E(n6453), .CP(clk), .QN(n18016) );
  EDFD1 \Mem_reg[59][30]  ( .D(n24783), .E(n6452), .CP(clk), .QN(n4972) );
  EDFD1 \Mem_reg[58][30]  ( .D(n24783), .E(n6451), .CP(clk), .QN(n4924) );
  EDFD1 \Mem_reg[57][30]  ( .D(n24783), .E(n6450), .CP(clk), .QN(n4876) );
  EDFD1 \Mem_reg[56][30]  ( .D(n24783), .E(n6449), .CP(clk), .QN(n4828) );
  EDFD1 \Mem_reg[55][30]  ( .D(n24783), .E(n6448), .CP(clk), .QN(n4780) );
  EDFD1 \Mem_reg[54][30]  ( .D(n24783), .E(n6447), .CP(clk), .QN(n15568) );
  EDFD1 \Mem_reg[53][30]  ( .D(n24783), .E(n6446), .CP(clk), .QN(n4684) );
  EDFD1 \Mem_reg[52][30]  ( .D(n24783), .E(n6445), .CP(clk), .Q(n27156) );
  EDFD1 \Mem_reg[51][30]  ( .D(n24783), .E(n6444), .CP(clk), .QN(n4588) );
  EDFD1 \Mem_reg[50][30]  ( .D(n24783), .E(n6443), .CP(clk), .QN(n4540) );
  EDFD1 \Mem_reg[49][30]  ( .D(n24783), .E(n6442), .CP(clk), .QN(n4492) );
  EDFD1 \Mem_reg[48][30]  ( .D(n24783), .E(n6441), .CP(clk), .QN(n4444) );
  EDFD1 \Mem_reg[47][30]  ( .D(n24783), .E(n6440), .CP(clk), .QN(n4396) );
  EDFD1 \Mem_reg[46][30]  ( .D(n24783), .E(n6439), .CP(clk), .QN(n4348) );
  EDFD1 \Mem_reg[43][30]  ( .D(n24783), .E(n6438), .CP(clk), .QN(n4300) );
  EDFD1 \Mem_reg[42][30]  ( .D(n24783), .E(n6437), .CP(clk), .QN(n4252) );
  EDFD1 \Mem_reg[41][30]  ( .D(n24783), .E(n6436), .CP(clk), .QN(n4204) );
  EDFD1 \Mem_reg[40][30]  ( .D(n24783), .E(n6435), .CP(clk), .QN(n4156) );
  EDFD1 \Mem_reg[39][30]  ( .D(n24783), .E(n6434), .CP(clk), .QN(n4108) );
  EDFD1 \Mem_reg[38][30]  ( .D(n24783), .E(n6433), .CP(clk), .QN(n4060) );
  EDFD1 \Mem_reg[37][30]  ( .D(n24783), .E(n6432), .CP(clk), .QN(n4012) );
  EDFD1 \Mem_reg[36][30]  ( .D(n24783), .E(n6431), .CP(clk), .QN(n3964) );
  EDFD1 \Mem_reg[35][30]  ( .D(n24783), .E(n6430), .CP(clk), .QN(n3916) );
  EDFD1 \Mem_reg[34][30]  ( .D(n24783), .E(n6429), .CP(clk), .QN(n3868) );
  EDFD1 \Mem_reg[33][30]  ( .D(n24783), .E(n6428), .CP(clk), .QN(n3820) );
  EDFD1 \Mem_reg[32][30]  ( .D(n24783), .E(n6427), .CP(clk), .QN(n3772) );
  EDFD1 \Mem_reg[31][30]  ( .D(n24783), .E(n6426), .CP(clk), .QN(n3724) );
  EDFD1 \Mem_reg[30][30]  ( .D(n24783), .E(n6425), .CP(clk), .QN(n3676) );
  EDFD1 \Mem_reg[29][30]  ( .D(n24783), .E(n6424), .CP(clk), .QN(n3628) );
  EDFD1 \Mem_reg[28][30]  ( .D(n24783), .E(n6423), .CP(clk), .QN(n3580) );
  EDFD1 \Mem_reg[27][30]  ( .D(n24783), .E(n6422), .CP(clk), .QN(n3532) );
  EDFD1 \Mem_reg[26][30]  ( .D(n24783), .E(n6421), .CP(clk), .QN(n3484) );
  EDFD1 \Mem_reg[25][30]  ( .D(n24783), .E(n6420), .CP(clk), .QN(n3436) );
  EDFD1 \Mem_reg[24][30]  ( .D(n24783), .E(n6463), .CP(clk), .QN(n3388) );
  EDFD1 \Mem_reg[23][30]  ( .D(n24783), .E(n6464), .CP(clk), .QN(n3340) );
  EDFD1 \Mem_reg[22][30]  ( .D(n24783), .E(n6465), .CP(clk), .QN(n3292) );
  EDFD1 \Mem_reg[21][30]  ( .D(n24783), .E(n6466), .CP(clk), .QN(n3244) );
  EDFD1 \Mem_reg[20][30]  ( .D(n24783), .E(n6467), .CP(clk), .QN(n3196) );
  EDFD1 \Mem_reg[19][30]  ( .D(n24783), .E(n6468), .CP(clk), .QN(n3148) );
  EDFD1 \Mem_reg[18][30]  ( .D(n24783), .E(n6469), .CP(clk), .QN(n3100) );
  EDFD1 \Mem_reg[17][30]  ( .D(n24783), .E(n6470), .CP(clk), .QN(n3052) );
  EDFD1 \Mem_reg[16][30]  ( .D(n24783), .E(n6471), .CP(clk), .QN(n3004) );
  EDFD1 \Mem_reg[15][30]  ( .D(n24783), .E(n6472), .CP(clk), .QN(n2956) );
  EDFD1 \Mem_reg[14][30]  ( .D(n24783), .E(n24720), .CP(clk), .QN(n2908) );
  EDFD1 \Mem_reg[13][30]  ( .D(n24783), .E(n24709), .CP(clk), .QN(n2860) );
  EDFD1 \Mem_reg[12][30]  ( .D(n24783), .E(n24717), .CP(clk), .QN(n2812) );
  EDFD1 \Mem_reg[11][30]  ( .D(n24783), .E(n24707), .CP(clk), .QN(n2764) );
  EDFD1 \Mem_reg[10][30]  ( .D(n24783), .E(n6477), .CP(clk), .QN(n2716) );
  EDFD1 \Mem_reg[9][30]  ( .D(n24783), .E(n24708), .CP(clk), .QN(n2668) );
  EDFD1 \Mem_reg[8][30]  ( .D(n24783), .E(n15642), .CP(clk), .QN(n2620) );
  EDFD1 \Mem_reg[7][30]  ( .D(n24783), .E(n24718), .CP(clk), .QN(n2572) );
  EDFD1 \Mem_reg[6][30]  ( .D(n24783), .E(n24716), .CP(clk), .QN(n2524) );
  EDFD1 \Mem_reg[5][30]  ( .D(n24783), .E(n24719), .CP(clk), .QN(n2476) );
  EDFD1 \Mem_reg[4][30]  ( .D(n24783), .E(n24706), .CP(clk), .QN(n2428) );
  EDFD1 \Mem_reg[3][30]  ( .D(n24783), .E(n24721), .CP(clk), .QN(n2380) );
  EDFD1 \Mem_reg[2][30]  ( .D(n24783), .E(n6460), .CP(clk), .QN(n2332) );
  EDFD1 \Mem_reg[1][30]  ( .D(n24783), .E(n24703), .CP(clk), .QN(n2284) );
  EDFD1 \Mem_reg[0][30]  ( .D(n24783), .E(n24705), .CP(clk), .QN(n2236) );
  EDFD1 \Mem_reg[88][29]  ( .D(n24781), .E(n6419), .CP(clk), .Q(n27153) );
  EDFD1 \Mem_reg[87][29]  ( .D(n24781), .E(n6418), .CP(clk), .QN(n6317) );
  EDFD1 \Mem_reg[86][29]  ( .D(n24781), .E(n6417), .CP(clk), .QN(n24646) );
  EDFD1 \Mem_reg[85][29]  ( .D(n24781), .E(n6416), .CP(clk), .QN(n6221) );
  EDFD1 \Mem_reg[84][29]  ( .D(n24781), .E(n6415), .CP(clk), .QN(n6173) );
  EDFD1 \Mem_reg[83][29]  ( .D(n24781), .E(n6414), .CP(clk), .QN(n6125) );
  EDFD1 \Mem_reg[82][29]  ( .D(n24781), .E(n6413), .CP(clk), .QN(n6077) );
  EDFD1 \Mem_reg[81][29]  ( .D(n24781), .E(n6412), .CP(clk), .QN(n6029) );
  EDFD1 \Mem_reg[80][29]  ( .D(n24781), .E(n6411), .CP(clk), .QN(n5981) );
  EDFD1 \Mem_reg[79][29]  ( .D(n24781), .E(n6410), .CP(clk), .QN(n5933) );
  EDFD1 \Mem_reg[78][29]  ( .D(n24781), .E(n6409), .CP(clk), .QN(n5885) );
  EDFD1 \Mem_reg[77][29]  ( .D(n24781), .E(n6408), .CP(clk), .QN(n5837) );
  EDFD1 \Mem_reg[76][29]  ( .D(n24781), .E(n6407), .CP(clk), .QN(n5789) );
  EDFD1 \Mem_reg[75][29]  ( .D(n24781), .E(n6406), .CP(clk), .QN(n27154) );
  EDFD1 \Mem_reg[74][29]  ( .D(n24781), .E(n6405), .CP(clk), .QN(n5693) );
  EDFD1 \Mem_reg[73][29]  ( .D(n24781), .E(n6404), .CP(clk), .QN(n27155) );
  EDFD1 \Mem_reg[72][29]  ( .D(n24781), .E(n6403), .CP(clk), .QN(n5597) );
  EDFD1 \Mem_reg[71][29]  ( .D(n24781), .E(n6402), .CP(clk), .QN(n5549) );
  EDFD1 \Mem_reg[70][29]  ( .D(n24781), .E(n6401), .CP(clk), .QN(n5501) );
  EDFD1 \Mem_reg[69][29]  ( .D(n24781), .E(n6400), .CP(clk), .QN(n5453) );
  EDFD1 \Mem_reg[68][29]  ( .D(n24781), .E(n6399), .CP(clk), .QN(n5405) );
  EDFD1 \Mem_reg[67][29]  ( .D(n24781), .E(n6398), .CP(clk), .QN(n5357) );
  EDFD1 \Mem_reg[66][29]  ( .D(n24781), .E(n6397), .CP(clk), .QN(n5309) );
  EDFD1 \Mem_reg[65][29]  ( .D(n24781), .E(n6396), .CP(clk), .QN(n15565) );
  EDFD1 \Mem_reg[64][29]  ( .D(n24781), .E(n6395), .CP(clk), .QN(n5213) );
  EDFD1 \Mem_reg[63][29]  ( .D(n24781), .E(n6456), .CP(clk), .QN(n5165) );
  EDFD1 \Mem_reg[62][29]  ( .D(n24781), .E(n6455), .CP(clk), .QN(n5117) );
  EDFD1 \Mem_reg[61][29]  ( .D(n24781), .E(n6454), .CP(clk), .QN(n18014) );
  EDFD1 \Mem_reg[60][29]  ( .D(n24781), .E(n6453), .CP(clk), .QN(n18013) );
  EDFD1 \Mem_reg[59][29]  ( .D(n24781), .E(n6452), .CP(clk), .QN(n4973) );
  EDFD1 \Mem_reg[58][29]  ( .D(n24781), .E(n6451), .CP(clk), .QN(n4925) );
  EDFD1 \Mem_reg[57][29]  ( .D(n24781), .E(n6450), .CP(clk), .QN(n4877) );
  EDFD1 \Mem_reg[56][29]  ( .D(n24781), .E(n6449), .CP(clk), .QN(n4829) );
  EDFD1 \Mem_reg[55][29]  ( .D(n24781), .E(n6448), .CP(clk), .QN(n4781) );
  EDFD1 \Mem_reg[54][29]  ( .D(n24781), .E(n6447), .CP(clk), .QN(n15564) );
  EDFD1 \Mem_reg[53][29]  ( .D(n24781), .E(n6446), .CP(clk), .QN(n4685) );
  EDFD1 \Mem_reg[52][29]  ( .D(n24781), .E(n6445), .CP(clk), .Q(n27152) );
  EDFD1 \Mem_reg[51][29]  ( .D(n24781), .E(n6444), .CP(clk), .QN(n4589) );
  EDFD1 \Mem_reg[50][29]  ( .D(n24781), .E(n6443), .CP(clk), .QN(n4541) );
  EDFD1 \Mem_reg[49][29]  ( .D(n24781), .E(n6442), .CP(clk), .QN(n4493) );
  EDFD1 \Mem_reg[48][29]  ( .D(n24781), .E(n6441), .CP(clk), .QN(n4445) );
  EDFD1 \Mem_reg[47][29]  ( .D(n24781), .E(n6440), .CP(clk), .QN(n4397) );
  EDFD1 \Mem_reg[46][29]  ( .D(n24781), .E(n6439), .CP(clk), .QN(n4349) );
  EDFD1 \Mem_reg[43][29]  ( .D(n24781), .E(n6438), .CP(clk), .QN(n4301) );
  EDFD1 \Mem_reg[42][29]  ( .D(n24781), .E(n6437), .CP(clk), .QN(n4253) );
  EDFD1 \Mem_reg[41][29]  ( .D(n24781), .E(n6436), .CP(clk), .QN(n4205) );
  EDFD1 \Mem_reg[40][29]  ( .D(n24781), .E(n6435), .CP(clk), .QN(n4157) );
  EDFD1 \Mem_reg[39][29]  ( .D(n24781), .E(n6434), .CP(clk), .QN(n4109) );
  EDFD1 \Mem_reg[38][29]  ( .D(n24781), .E(n6433), .CP(clk), .QN(n4061) );
  EDFD1 \Mem_reg[37][29]  ( .D(n24781), .E(n6432), .CP(clk), .QN(n4013) );
  EDFD1 \Mem_reg[36][29]  ( .D(n24781), .E(n6431), .CP(clk), .QN(n3965) );
  EDFD1 \Mem_reg[35][29]  ( .D(n24781), .E(n6430), .CP(clk), .QN(n3917) );
  EDFD1 \Mem_reg[34][29]  ( .D(n24781), .E(n6429), .CP(clk), .QN(n3869) );
  EDFD1 \Mem_reg[33][29]  ( .D(n24781), .E(n6428), .CP(clk), .QN(n3821) );
  EDFD1 \Mem_reg[32][29]  ( .D(n24781), .E(n6427), .CP(clk), .QN(n3773) );
  EDFD1 \Mem_reg[31][29]  ( .D(n24781), .E(n6426), .CP(clk), .QN(n3725) );
  EDFD1 \Mem_reg[30][29]  ( .D(n24781), .E(n6425), .CP(clk), .QN(n3677) );
  EDFD1 \Mem_reg[29][29]  ( .D(n24781), .E(n6424), .CP(clk), .QN(n3629) );
  EDFD1 \Mem_reg[28][29]  ( .D(n24781), .E(n6423), .CP(clk), .QN(n3581) );
  EDFD1 \Mem_reg[27][29]  ( .D(n24781), .E(n6422), .CP(clk), .QN(n3533) );
  EDFD1 \Mem_reg[26][29]  ( .D(n24781), .E(n6421), .CP(clk), .QN(n3485) );
  EDFD1 \Mem_reg[25][29]  ( .D(n24781), .E(n6420), .CP(clk), .QN(n3437) );
  EDFD1 \Mem_reg[24][29]  ( .D(n24781), .E(n6463), .CP(clk), .QN(n3389) );
  EDFD1 \Mem_reg[23][29]  ( .D(n24781), .E(n6464), .CP(clk), .QN(n3341) );
  EDFD1 \Mem_reg[22][29]  ( .D(n24781), .E(n6465), .CP(clk), .QN(n3293) );
  EDFD1 \Mem_reg[21][29]  ( .D(n24781), .E(n6466), .CP(clk), .QN(n3245) );
  EDFD1 \Mem_reg[20][29]  ( .D(n24781), .E(n6467), .CP(clk), .QN(n3197) );
  EDFD1 \Mem_reg[19][29]  ( .D(n24781), .E(n6468), .CP(clk), .QN(n3149) );
  EDFD1 \Mem_reg[18][29]  ( .D(n24781), .E(n6469), .CP(clk), .QN(n3101) );
  EDFD1 \Mem_reg[17][29]  ( .D(n24781), .E(n6470), .CP(clk), .QN(n3053) );
  EDFD1 \Mem_reg[16][29]  ( .D(n24781), .E(n6471), .CP(clk), .QN(n3005) );
  EDFD1 \Mem_reg[15][29]  ( .D(n24781), .E(n6472), .CP(clk), .QN(n2957) );
  EDFD1 \Mem_reg[14][29]  ( .D(n24781), .E(n24720), .CP(clk), .QN(n2909) );
  EDFD1 \Mem_reg[13][29]  ( .D(n24781), .E(n24709), .CP(clk), .QN(n2861) );
  EDFD1 \Mem_reg[12][29]  ( .D(n24781), .E(n24717), .CP(clk), .QN(n2813) );
  EDFD1 \Mem_reg[11][29]  ( .D(n24781), .E(n24707), .CP(clk), .QN(n2765) );
  EDFD1 \Mem_reg[10][29]  ( .D(n24781), .E(n6477), .CP(clk), .QN(n2717) );
  EDFD1 \Mem_reg[9][29]  ( .D(n24781), .E(n24708), .CP(clk), .QN(n2669) );
  EDFD1 \Mem_reg[8][29]  ( .D(n24781), .E(n15642), .CP(clk), .QN(n2621) );
  EDFD1 \Mem_reg[7][29]  ( .D(n24781), .E(n24718), .CP(clk), .QN(n2573) );
  EDFD1 \Mem_reg[6][29]  ( .D(n24781), .E(n24716), .CP(clk), .QN(n2525) );
  EDFD1 \Mem_reg[5][29]  ( .D(n24781), .E(n24719), .CP(clk), .QN(n2477) );
  EDFD1 \Mem_reg[4][29]  ( .D(n24781), .E(n24706), .CP(clk), .QN(n2429) );
  EDFD1 \Mem_reg[3][29]  ( .D(n24781), .E(n24721), .CP(clk), .QN(n2381) );
  EDFD1 \Mem_reg[2][29]  ( .D(n24781), .E(n6460), .CP(clk), .QN(n2333) );
  EDFD1 \Mem_reg[1][29]  ( .D(n24781), .E(n24703), .CP(clk), .QN(n2285) );
  EDFD1 \Mem_reg[0][29]  ( .D(n24781), .E(n24705), .CP(clk), .QN(n2237) );
  EDFD1 \Mem_reg[88][28]  ( .D(n24779), .E(n6419), .CP(clk), .Q(n27149) );
  EDFD1 \Mem_reg[87][28]  ( .D(n24779), .E(n6418), .CP(clk), .QN(n6318) );
  EDFD1 \Mem_reg[86][28]  ( .D(n24779), .E(n6417), .CP(clk), .QN(n24643) );
  EDFD1 \Mem_reg[85][28]  ( .D(n24779), .E(n6416), .CP(clk), .QN(n6222) );
  EDFD1 \Mem_reg[84][28]  ( .D(n24779), .E(n6415), .CP(clk), .QN(n6174) );
  EDFD1 \Mem_reg[83][28]  ( .D(n24779), .E(n6414), .CP(clk), .QN(n6126) );
  EDFD1 \Mem_reg[82][28]  ( .D(n24779), .E(n6413), .CP(clk), .QN(n6078) );
  EDFD1 \Mem_reg[81][28]  ( .D(n24779), .E(n6412), .CP(clk), .QN(n6030) );
  EDFD1 \Mem_reg[80][28]  ( .D(n24779), .E(n6411), .CP(clk), .QN(n5982) );
  EDFD1 \Mem_reg[79][28]  ( .D(n24779), .E(n6410), .CP(clk), .QN(n5934) );
  EDFD1 \Mem_reg[78][28]  ( .D(n24779), .E(n6409), .CP(clk), .QN(n5886) );
  EDFD1 \Mem_reg[77][28]  ( .D(n24779), .E(n6408), .CP(clk), .QN(n5838) );
  EDFD1 \Mem_reg[76][28]  ( .D(n24779), .E(n6407), .CP(clk), .QN(n5790) );
  EDFD1 \Mem_reg[75][28]  ( .D(n24779), .E(n6406), .CP(clk), .QN(n27150) );
  EDFD1 \Mem_reg[74][28]  ( .D(n24779), .E(n6405), .CP(clk), .QN(n5694) );
  EDFD1 \Mem_reg[73][28]  ( .D(n24779), .E(n6404), .CP(clk), .QN(n27151) );
  EDFD1 \Mem_reg[72][28]  ( .D(n24779), .E(n6403), .CP(clk), .QN(n5598) );
  EDFD1 \Mem_reg[71][28]  ( .D(n24779), .E(n6402), .CP(clk), .QN(n5550) );
  EDFD1 \Mem_reg[70][28]  ( .D(n24779), .E(n6401), .CP(clk), .QN(n5502) );
  EDFD1 \Mem_reg[69][28]  ( .D(n24779), .E(n6400), .CP(clk), .QN(n5454) );
  EDFD1 \Mem_reg[68][28]  ( .D(n24779), .E(n6399), .CP(clk), .QN(n5406) );
  EDFD1 \Mem_reg[67][28]  ( .D(n24779), .E(n6398), .CP(clk), .QN(n5358) );
  EDFD1 \Mem_reg[66][28]  ( .D(n24779), .E(n6397), .CP(clk), .QN(n5310) );
  EDFD1 \Mem_reg[65][28]  ( .D(n24779), .E(n6396), .CP(clk), .QN(n15561) );
  EDFD1 \Mem_reg[64][28]  ( .D(n24779), .E(n6395), .CP(clk), .QN(n5214) );
  EDFD1 \Mem_reg[63][28]  ( .D(n24779), .E(n6456), .CP(clk), .QN(n5166) );
  EDFD1 \Mem_reg[62][28]  ( .D(n24779), .E(n6455), .CP(clk), .QN(n5118) );
  EDFD1 \Mem_reg[61][28]  ( .D(n24779), .E(n6454), .CP(clk), .QN(n18011) );
  EDFD1 \Mem_reg[60][28]  ( .D(n24779), .E(n6453), .CP(clk), .QN(n18010) );
  EDFD1 \Mem_reg[59][28]  ( .D(n24779), .E(n6452), .CP(clk), .QN(n4974) );
  EDFD1 \Mem_reg[58][28]  ( .D(n24779), .E(n6451), .CP(clk), .QN(n4926) );
  EDFD1 \Mem_reg[57][28]  ( .D(n24779), .E(n6450), .CP(clk), .QN(n4878) );
  EDFD1 \Mem_reg[56][28]  ( .D(n24779), .E(n6449), .CP(clk), .QN(n4830) );
  EDFD1 \Mem_reg[55][28]  ( .D(n24779), .E(n6448), .CP(clk), .QN(n4782) );
  EDFD1 \Mem_reg[54][28]  ( .D(n24779), .E(n6447), .CP(clk), .QN(n15560) );
  EDFD1 \Mem_reg[53][28]  ( .D(n24779), .E(n6446), .CP(clk), .QN(n4686) );
  EDFD1 \Mem_reg[52][28]  ( .D(n24779), .E(n6445), .CP(clk), .Q(n27148) );
  EDFD1 \Mem_reg[51][28]  ( .D(n24779), .E(n6444), .CP(clk), .QN(n4590) );
  EDFD1 \Mem_reg[50][28]  ( .D(n24779), .E(n6443), .CP(clk), .QN(n4542) );
  EDFD1 \Mem_reg[49][28]  ( .D(n24779), .E(n6442), .CP(clk), .QN(n4494) );
  EDFD1 \Mem_reg[48][28]  ( .D(n24779), .E(n6441), .CP(clk), .QN(n4446) );
  EDFD1 \Mem_reg[47][28]  ( .D(n24779), .E(n6440), .CP(clk), .QN(n4398) );
  EDFD1 \Mem_reg[46][28]  ( .D(n24779), .E(n6439), .CP(clk), .QN(n4350) );
  EDFD1 \Mem_reg[43][28]  ( .D(n24779), .E(n6438), .CP(clk), .QN(n4302) );
  EDFD1 \Mem_reg[42][28]  ( .D(n24779), .E(n6437), .CP(clk), .QN(n4254) );
  EDFD1 \Mem_reg[41][28]  ( .D(n24779), .E(n6436), .CP(clk), .QN(n4206) );
  EDFD1 \Mem_reg[40][28]  ( .D(n24779), .E(n6435), .CP(clk), .QN(n4158) );
  EDFD1 \Mem_reg[39][28]  ( .D(n24779), .E(n6434), .CP(clk), .QN(n4110) );
  EDFD1 \Mem_reg[38][28]  ( .D(n24779), .E(n6433), .CP(clk), .QN(n4062) );
  EDFD1 \Mem_reg[37][28]  ( .D(n24779), .E(n6432), .CP(clk), .QN(n4014) );
  EDFD1 \Mem_reg[36][28]  ( .D(n24779), .E(n6431), .CP(clk), .QN(n3966) );
  EDFD1 \Mem_reg[35][28]  ( .D(n24779), .E(n6430), .CP(clk), .QN(n3918) );
  EDFD1 \Mem_reg[34][28]  ( .D(n24779), .E(n6429), .CP(clk), .QN(n3870) );
  EDFD1 \Mem_reg[33][28]  ( .D(n24779), .E(n6428), .CP(clk), .QN(n3822) );
  EDFD1 \Mem_reg[32][28]  ( .D(n24779), .E(n6427), .CP(clk), .QN(n3774) );
  EDFD1 \Mem_reg[31][28]  ( .D(n24779), .E(n6426), .CP(clk), .QN(n3726) );
  EDFD1 \Mem_reg[30][28]  ( .D(n24779), .E(n6425), .CP(clk), .QN(n3678) );
  EDFD1 \Mem_reg[29][28]  ( .D(n24779), .E(n6424), .CP(clk), .QN(n3630) );
  EDFD1 \Mem_reg[28][28]  ( .D(n24779), .E(n6423), .CP(clk), .QN(n3582) );
  EDFD1 \Mem_reg[27][28]  ( .D(n24779), .E(n6422), .CP(clk), .QN(n3534) );
  EDFD1 \Mem_reg[26][28]  ( .D(n24779), .E(n6421), .CP(clk), .QN(n3486) );
  EDFD1 \Mem_reg[25][28]  ( .D(n24779), .E(n6420), .CP(clk), .QN(n3438) );
  EDFD1 \Mem_reg[24][28]  ( .D(n24779), .E(n6463), .CP(clk), .QN(n3390) );
  EDFD1 \Mem_reg[23][28]  ( .D(n24779), .E(n6464), .CP(clk), .QN(n3342) );
  EDFD1 \Mem_reg[22][28]  ( .D(n24779), .E(n6465), .CP(clk), .QN(n3294) );
  EDFD1 \Mem_reg[21][28]  ( .D(n24779), .E(n6466), .CP(clk), .QN(n3246) );
  EDFD1 \Mem_reg[20][28]  ( .D(n24779), .E(n6467), .CP(clk), .QN(n3198) );
  EDFD1 \Mem_reg[19][28]  ( .D(n24779), .E(n6468), .CP(clk), .QN(n3150) );
  EDFD1 \Mem_reg[18][28]  ( .D(n24779), .E(n6469), .CP(clk), .QN(n3102) );
  EDFD1 \Mem_reg[17][28]  ( .D(n24779), .E(n6470), .CP(clk), .QN(n3054) );
  EDFD1 \Mem_reg[16][28]  ( .D(n24779), .E(n6471), .CP(clk), .QN(n3006) );
  EDFD1 \Mem_reg[15][28]  ( .D(n24779), .E(n6472), .CP(clk), .QN(n2958) );
  EDFD1 \Mem_reg[14][28]  ( .D(n24779), .E(n24720), .CP(clk), .QN(n2910) );
  EDFD1 \Mem_reg[13][28]  ( .D(n24779), .E(n24709), .CP(clk), .QN(n2862) );
  EDFD1 \Mem_reg[12][28]  ( .D(n24779), .E(n24717), .CP(clk), .QN(n2814) );
  EDFD1 \Mem_reg[11][28]  ( .D(n24779), .E(n24707), .CP(clk), .QN(n2766) );
  EDFD1 \Mem_reg[10][28]  ( .D(n24779), .E(n6477), .CP(clk), .QN(n2718) );
  EDFD1 \Mem_reg[9][28]  ( .D(n24779), .E(n24708), .CP(clk), .QN(n2670) );
  EDFD1 \Mem_reg[8][28]  ( .D(n24779), .E(n15642), .CP(clk), .QN(n2622) );
  EDFD1 \Mem_reg[7][28]  ( .D(n24779), .E(n24718), .CP(clk), .QN(n2574) );
  EDFD1 \Mem_reg[6][28]  ( .D(n24779), .E(n24716), .CP(clk), .QN(n2526) );
  EDFD1 \Mem_reg[5][28]  ( .D(n24779), .E(n24719), .CP(clk), .QN(n2478) );
  EDFD1 \Mem_reg[4][28]  ( .D(n24779), .E(n24706), .CP(clk), .QN(n2430) );
  EDFD1 \Mem_reg[3][28]  ( .D(n24779), .E(n24721), .CP(clk), .QN(n2382) );
  EDFD1 \Mem_reg[2][28]  ( .D(n24779), .E(n6460), .CP(clk), .QN(n2334) );
  EDFD1 \Mem_reg[1][28]  ( .D(n24779), .E(n24703), .CP(clk), .QN(n2286) );
  EDFD1 \Mem_reg[0][28]  ( .D(n24779), .E(n24705), .CP(clk), .QN(n2238) );
  EDFD1 \Mem_reg[88][27]  ( .D(n24777), .E(n6419), .CP(clk), .Q(n27145) );
  EDFD1 \Mem_reg[87][27]  ( .D(n24777), .E(n6418), .CP(clk), .QN(n6319) );
  EDFD1 \Mem_reg[86][27]  ( .D(n24777), .E(n6417), .CP(clk), .QN(n24640) );
  EDFD1 \Mem_reg[85][27]  ( .D(n24777), .E(n6416), .CP(clk), .QN(n6223) );
  EDFD1 \Mem_reg[84][27]  ( .D(n24777), .E(n6415), .CP(clk), .QN(n6175) );
  EDFD1 \Mem_reg[83][27]  ( .D(n24777), .E(n6414), .CP(clk), .QN(n6127) );
  EDFD1 \Mem_reg[82][27]  ( .D(n24777), .E(n6413), .CP(clk), .QN(n6079) );
  EDFD1 \Mem_reg[81][27]  ( .D(n24777), .E(n6412), .CP(clk), .QN(n6031) );
  EDFD1 \Mem_reg[80][27]  ( .D(n24777), .E(n6411), .CP(clk), .QN(n5983) );
  EDFD1 \Mem_reg[79][27]  ( .D(n24777), .E(n6410), .CP(clk), .QN(n5935) );
  EDFD1 \Mem_reg[78][27]  ( .D(n24777), .E(n6409), .CP(clk), .QN(n5887) );
  EDFD1 \Mem_reg[77][27]  ( .D(n24777), .E(n6408), .CP(clk), .QN(n5839) );
  EDFD1 \Mem_reg[76][27]  ( .D(n24777), .E(n6407), .CP(clk), .QN(n5791) );
  EDFD1 \Mem_reg[75][27]  ( .D(n24777), .E(n6406), .CP(clk), .QN(n27146) );
  EDFD1 \Mem_reg[74][27]  ( .D(n24777), .E(n6405), .CP(clk), .QN(n5695) );
  EDFD1 \Mem_reg[73][27]  ( .D(n24777), .E(n6404), .CP(clk), .QN(n27147) );
  EDFD1 \Mem_reg[72][27]  ( .D(n24777), .E(n6403), .CP(clk), .QN(n5599) );
  EDFD1 \Mem_reg[71][27]  ( .D(n24777), .E(n6402), .CP(clk), .QN(n5551) );
  EDFD1 \Mem_reg[70][27]  ( .D(n24777), .E(n6401), .CP(clk), .QN(n5503) );
  EDFD1 \Mem_reg[69][27]  ( .D(n24777), .E(n6400), .CP(clk), .QN(n5455) );
  EDFD1 \Mem_reg[68][27]  ( .D(n24777), .E(n6399), .CP(clk), .QN(n5407) );
  EDFD1 \Mem_reg[67][27]  ( .D(n24777), .E(n6398), .CP(clk), .QN(n5359) );
  EDFD1 \Mem_reg[66][27]  ( .D(n24777), .E(n6397), .CP(clk), .QN(n5311) );
  EDFD1 \Mem_reg[65][27]  ( .D(n24777), .E(n6396), .CP(clk), .QN(n15557) );
  EDFD1 \Mem_reg[64][27]  ( .D(n24777), .E(n6395), .CP(clk), .QN(n5215) );
  EDFD1 \Mem_reg[63][27]  ( .D(n24777), .E(n6456), .CP(clk), .QN(n5167) );
  EDFD1 \Mem_reg[62][27]  ( .D(n24777), .E(n6455), .CP(clk), .QN(n5119) );
  EDFD1 \Mem_reg[61][27]  ( .D(n24777), .E(n6454), .CP(clk), .QN(n18008) );
  EDFD1 \Mem_reg[60][27]  ( .D(n24777), .E(n6453), .CP(clk), .QN(n18007) );
  EDFD1 \Mem_reg[59][27]  ( .D(n24777), .E(n6452), .CP(clk), .QN(n4975) );
  EDFD1 \Mem_reg[58][27]  ( .D(n24777), .E(n6451), .CP(clk), .QN(n4927) );
  EDFD1 \Mem_reg[57][27]  ( .D(n24777), .E(n6450), .CP(clk), .QN(n4879) );
  EDFD1 \Mem_reg[56][27]  ( .D(n24777), .E(n6449), .CP(clk), .QN(n4831) );
  EDFD1 \Mem_reg[55][27]  ( .D(n24777), .E(n6448), .CP(clk), .QN(n4783) );
  EDFD1 \Mem_reg[54][27]  ( .D(n24777), .E(n6447), .CP(clk), .QN(n15556) );
  EDFD1 \Mem_reg[53][27]  ( .D(n24777), .E(n6446), .CP(clk), .QN(n4687) );
  EDFD1 \Mem_reg[52][27]  ( .D(n24777), .E(n6445), .CP(clk), .Q(n27144) );
  EDFD1 \Mem_reg[51][27]  ( .D(n24777), .E(n6444), .CP(clk), .QN(n4591) );
  EDFD1 \Mem_reg[50][27]  ( .D(n24777), .E(n6443), .CP(clk), .QN(n4543) );
  EDFD1 \Mem_reg[49][27]  ( .D(n24777), .E(n6442), .CP(clk), .QN(n4495) );
  EDFD1 \Mem_reg[48][27]  ( .D(n24777), .E(n6441), .CP(clk), .QN(n4447) );
  EDFD1 \Mem_reg[47][27]  ( .D(n24777), .E(n6440), .CP(clk), .QN(n4399) );
  EDFD1 \Mem_reg[46][27]  ( .D(n24777), .E(n6439), .CP(clk), .QN(n4351) );
  EDFD1 \Mem_reg[43][27]  ( .D(n24777), .E(n6438), .CP(clk), .QN(n4303) );
  EDFD1 \Mem_reg[42][27]  ( .D(n24777), .E(n6437), .CP(clk), .QN(n4255) );
  EDFD1 \Mem_reg[41][27]  ( .D(n24777), .E(n6436), .CP(clk), .QN(n4207) );
  EDFD1 \Mem_reg[40][27]  ( .D(n24777), .E(n6435), .CP(clk), .QN(n4159) );
  EDFD1 \Mem_reg[39][27]  ( .D(n24777), .E(n6434), .CP(clk), .QN(n4111) );
  EDFD1 \Mem_reg[38][27]  ( .D(n24777), .E(n6433), .CP(clk), .QN(n4063) );
  EDFD1 \Mem_reg[37][27]  ( .D(n24777), .E(n6432), .CP(clk), .QN(n4015) );
  EDFD1 \Mem_reg[36][27]  ( .D(n24777), .E(n6431), .CP(clk), .QN(n3967) );
  EDFD1 \Mem_reg[35][27]  ( .D(n24777), .E(n6430), .CP(clk), .QN(n3919) );
  EDFD1 \Mem_reg[34][27]  ( .D(n24777), .E(n6429), .CP(clk), .QN(n3871) );
  EDFD1 \Mem_reg[33][27]  ( .D(n24777), .E(n6428), .CP(clk), .QN(n3823) );
  EDFD1 \Mem_reg[32][27]  ( .D(n24777), .E(n6427), .CP(clk), .QN(n3775) );
  EDFD1 \Mem_reg[31][27]  ( .D(n24777), .E(n6426), .CP(clk), .QN(n3727) );
  EDFD1 \Mem_reg[30][27]  ( .D(n24777), .E(n6425), .CP(clk), .QN(n3679) );
  EDFD1 \Mem_reg[29][27]  ( .D(n24777), .E(n6424), .CP(clk), .QN(n3631) );
  EDFD1 \Mem_reg[28][27]  ( .D(n24777), .E(n6423), .CP(clk), .QN(n3583) );
  EDFD1 \Mem_reg[27][27]  ( .D(n24777), .E(n6422), .CP(clk), .QN(n3535) );
  EDFD1 \Mem_reg[26][27]  ( .D(n24777), .E(n6421), .CP(clk), .QN(n3487) );
  EDFD1 \Mem_reg[25][27]  ( .D(n24777), .E(n6420), .CP(clk), .QN(n3439) );
  EDFD1 \Mem_reg[24][27]  ( .D(n24777), .E(n6463), .CP(clk), .QN(n3391) );
  EDFD1 \Mem_reg[23][27]  ( .D(n24777), .E(n6464), .CP(clk), .QN(n3343) );
  EDFD1 \Mem_reg[22][27]  ( .D(n24777), .E(n6465), .CP(clk), .QN(n3295) );
  EDFD1 \Mem_reg[21][27]  ( .D(n24777), .E(n6466), .CP(clk), .QN(n3247) );
  EDFD1 \Mem_reg[20][27]  ( .D(n24777), .E(n6467), .CP(clk), .QN(n3199) );
  EDFD1 \Mem_reg[19][27]  ( .D(n24777), .E(n6468), .CP(clk), .QN(n3151) );
  EDFD1 \Mem_reg[18][27]  ( .D(n24777), .E(n6469), .CP(clk), .QN(n3103) );
  EDFD1 \Mem_reg[17][27]  ( .D(n24777), .E(n6470), .CP(clk), .QN(n3055) );
  EDFD1 \Mem_reg[16][27]  ( .D(n24777), .E(n6471), .CP(clk), .QN(n3007) );
  EDFD1 \Mem_reg[15][27]  ( .D(n24777), .E(n6472), .CP(clk), .QN(n2959) );
  EDFD1 \Mem_reg[14][27]  ( .D(n24777), .E(n24720), .CP(clk), .QN(n2911) );
  EDFD1 \Mem_reg[13][27]  ( .D(n24777), .E(n24709), .CP(clk), .QN(n2863) );
  EDFD1 \Mem_reg[12][27]  ( .D(n24777), .E(n24717), .CP(clk), .QN(n2815) );
  EDFD1 \Mem_reg[11][27]  ( .D(n24777), .E(n24707), .CP(clk), .QN(n2767) );
  EDFD1 \Mem_reg[10][27]  ( .D(n24777), .E(n6477), .CP(clk), .QN(n2719) );
  EDFD1 \Mem_reg[9][27]  ( .D(n24777), .E(n24708), .CP(clk), .QN(n2671) );
  EDFD1 \Mem_reg[8][27]  ( .D(n24777), .E(n15642), .CP(clk), .QN(n2623) );
  EDFD1 \Mem_reg[7][27]  ( .D(n24777), .E(n24718), .CP(clk), .QN(n2575) );
  EDFD1 \Mem_reg[6][27]  ( .D(n24777), .E(n24716), .CP(clk), .QN(n2527) );
  EDFD1 \Mem_reg[5][27]  ( .D(n24777), .E(n24719), .CP(clk), .QN(n2479) );
  EDFD1 \Mem_reg[4][27]  ( .D(n24777), .E(n24706), .CP(clk), .QN(n2431) );
  EDFD1 \Mem_reg[3][27]  ( .D(n24777), .E(n24721), .CP(clk), .QN(n2383) );
  EDFD1 \Mem_reg[2][27]  ( .D(n24777), .E(n6460), .CP(clk), .QN(n2335) );
  EDFD1 \Mem_reg[1][27]  ( .D(n24777), .E(n24703), .CP(clk), .QN(n2287) );
  EDFD1 \Mem_reg[0][27]  ( .D(n24777), .E(n24705), .CP(clk), .QN(n2239) );
  EDFD1 \Mem_reg[88][26]  ( .D(n24775), .E(n6419), .CP(clk), .Q(n27141) );
  EDFD1 \Mem_reg[87][26]  ( .D(n24775), .E(n6418), .CP(clk), .QN(n6320) );
  EDFD1 \Mem_reg[86][26]  ( .D(n24775), .E(n6417), .CP(clk), .QN(n24637) );
  EDFD1 \Mem_reg[85][26]  ( .D(n24775), .E(n6416), .CP(clk), .QN(n6224) );
  EDFD1 \Mem_reg[84][26]  ( .D(n24775), .E(n6415), .CP(clk), .QN(n6176) );
  EDFD1 \Mem_reg[83][26]  ( .D(n24775), .E(n6414), .CP(clk), .QN(n6128) );
  EDFD1 \Mem_reg[82][26]  ( .D(n24775), .E(n6413), .CP(clk), .QN(n6080) );
  EDFD1 \Mem_reg[81][26]  ( .D(n24775), .E(n6412), .CP(clk), .QN(n6032) );
  EDFD1 \Mem_reg[80][26]  ( .D(n24775), .E(n6411), .CP(clk), .QN(n5984) );
  EDFD1 \Mem_reg[79][26]  ( .D(n24775), .E(n6410), .CP(clk), .QN(n5936) );
  EDFD1 \Mem_reg[78][26]  ( .D(n24775), .E(n6409), .CP(clk), .QN(n5888) );
  EDFD1 \Mem_reg[77][26]  ( .D(n24775), .E(n6408), .CP(clk), .QN(n5840) );
  EDFD1 \Mem_reg[76][26]  ( .D(n24775), .E(n6407), .CP(clk), .QN(n5792) );
  EDFD1 \Mem_reg[75][26]  ( .D(n24775), .E(n6406), .CP(clk), .QN(n27142) );
  EDFD1 \Mem_reg[74][26]  ( .D(n24775), .E(n6405), .CP(clk), .QN(n5696) );
  EDFD1 \Mem_reg[73][26]  ( .D(n24775), .E(n6404), .CP(clk), .QN(n27143) );
  EDFD1 \Mem_reg[72][26]  ( .D(n24775), .E(n6403), .CP(clk), .QN(n5600) );
  EDFD1 \Mem_reg[71][26]  ( .D(n24775), .E(n6402), .CP(clk), .QN(n5552) );
  EDFD1 \Mem_reg[70][26]  ( .D(n24775), .E(n6401), .CP(clk), .QN(n5504) );
  EDFD1 \Mem_reg[69][26]  ( .D(n24775), .E(n6400), .CP(clk), .QN(n5456) );
  EDFD1 \Mem_reg[68][26]  ( .D(n24775), .E(n6399), .CP(clk), .QN(n5408) );
  EDFD1 \Mem_reg[67][26]  ( .D(n24775), .E(n6398), .CP(clk), .QN(n5360) );
  EDFD1 \Mem_reg[66][26]  ( .D(n24775), .E(n6397), .CP(clk), .QN(n5312) );
  EDFD1 \Mem_reg[65][26]  ( .D(n24775), .E(n6396), .CP(clk), .QN(n15553) );
  EDFD1 \Mem_reg[64][26]  ( .D(n24775), .E(n6395), .CP(clk), .QN(n5216) );
  EDFD1 \Mem_reg[63][26]  ( .D(n24775), .E(n6456), .CP(clk), .QN(n5168) );
  EDFD1 \Mem_reg[62][26]  ( .D(n24775), .E(n6455), .CP(clk), .QN(n5120) );
  EDFD1 \Mem_reg[61][26]  ( .D(n24775), .E(n6454), .CP(clk), .QN(n18005) );
  EDFD1 \Mem_reg[60][26]  ( .D(n24775), .E(n6453), .CP(clk), .QN(n18004) );
  EDFD1 \Mem_reg[59][26]  ( .D(n24775), .E(n6452), .CP(clk), .QN(n4976) );
  EDFD1 \Mem_reg[58][26]  ( .D(n24775), .E(n6451), .CP(clk), .QN(n4928) );
  EDFD1 \Mem_reg[57][26]  ( .D(n24775), .E(n6450), .CP(clk), .QN(n4880) );
  EDFD1 \Mem_reg[56][26]  ( .D(n24775), .E(n6449), .CP(clk), .QN(n4832) );
  EDFD1 \Mem_reg[55][26]  ( .D(n24775), .E(n6448), .CP(clk), .QN(n4784) );
  EDFD1 \Mem_reg[54][26]  ( .D(n24775), .E(n6447), .CP(clk), .QN(n15552) );
  EDFD1 \Mem_reg[53][26]  ( .D(n24775), .E(n6446), .CP(clk), .QN(n4688) );
  EDFD1 \Mem_reg[52][26]  ( .D(n24775), .E(n6445), .CP(clk), .Q(n27140) );
  EDFD1 \Mem_reg[51][26]  ( .D(n24775), .E(n6444), .CP(clk), .QN(n4592) );
  EDFD1 \Mem_reg[50][26]  ( .D(n24775), .E(n6443), .CP(clk), .QN(n4544) );
  EDFD1 \Mem_reg[49][26]  ( .D(n24775), .E(n6442), .CP(clk), .QN(n4496) );
  EDFD1 \Mem_reg[48][26]  ( .D(n24775), .E(n6441), .CP(clk), .QN(n4448) );
  EDFD1 \Mem_reg[47][26]  ( .D(n24775), .E(n6440), .CP(clk), .QN(n4400) );
  EDFD1 \Mem_reg[46][26]  ( .D(n24775), .E(n6439), .CP(clk), .QN(n4352) );
  EDFD1 \Mem_reg[43][26]  ( .D(n24775), .E(n6438), .CP(clk), .QN(n4304) );
  EDFD1 \Mem_reg[42][26]  ( .D(n24775), .E(n6437), .CP(clk), .QN(n4256) );
  EDFD1 \Mem_reg[41][26]  ( .D(n24775), .E(n6436), .CP(clk), .QN(n4208) );
  EDFD1 \Mem_reg[40][26]  ( .D(n24775), .E(n6435), .CP(clk), .QN(n4160) );
  EDFD1 \Mem_reg[39][26]  ( .D(n24775), .E(n6434), .CP(clk), .QN(n4112) );
  EDFD1 \Mem_reg[38][26]  ( .D(n24775), .E(n6433), .CP(clk), .QN(n4064) );
  EDFD1 \Mem_reg[37][26]  ( .D(n24775), .E(n6432), .CP(clk), .QN(n4016) );
  EDFD1 \Mem_reg[36][26]  ( .D(n24775), .E(n6431), .CP(clk), .QN(n3968) );
  EDFD1 \Mem_reg[35][26]  ( .D(n24775), .E(n6430), .CP(clk), .QN(n3920) );
  EDFD1 \Mem_reg[34][26]  ( .D(n24775), .E(n6429), .CP(clk), .QN(n3872) );
  EDFD1 \Mem_reg[33][26]  ( .D(n24775), .E(n6428), .CP(clk), .QN(n3824) );
  EDFD1 \Mem_reg[32][26]  ( .D(n24775), .E(n6427), .CP(clk), .QN(n3776) );
  EDFD1 \Mem_reg[31][26]  ( .D(n24775), .E(n6426), .CP(clk), .QN(n3728) );
  EDFD1 \Mem_reg[30][26]  ( .D(n24775), .E(n6425), .CP(clk), .QN(n3680) );
  EDFD1 \Mem_reg[29][26]  ( .D(n24775), .E(n6424), .CP(clk), .QN(n3632) );
  EDFD1 \Mem_reg[28][26]  ( .D(n24775), .E(n6423), .CP(clk), .QN(n3584) );
  EDFD1 \Mem_reg[27][26]  ( .D(n24775), .E(n6422), .CP(clk), .QN(n3536) );
  EDFD1 \Mem_reg[26][26]  ( .D(n24775), .E(n6421), .CP(clk), .QN(n3488) );
  EDFD1 \Mem_reg[25][26]  ( .D(n24775), .E(n6420), .CP(clk), .QN(n3440) );
  EDFD1 \Mem_reg[24][26]  ( .D(n24775), .E(n6463), .CP(clk), .QN(n3392) );
  EDFD1 \Mem_reg[23][26]  ( .D(n24775), .E(n6464), .CP(clk), .QN(n3344) );
  EDFD1 \Mem_reg[22][26]  ( .D(n24775), .E(n6465), .CP(clk), .QN(n3296) );
  EDFD1 \Mem_reg[21][26]  ( .D(n24775), .E(n6466), .CP(clk), .QN(n3248) );
  EDFD1 \Mem_reg[20][26]  ( .D(n24775), .E(n6467), .CP(clk), .QN(n3200) );
  EDFD1 \Mem_reg[19][26]  ( .D(n24775), .E(n6468), .CP(clk), .QN(n3152) );
  EDFD1 \Mem_reg[18][26]  ( .D(n24775), .E(n6469), .CP(clk), .QN(n3104) );
  EDFD1 \Mem_reg[17][26]  ( .D(n24775), .E(n6470), .CP(clk), .QN(n3056) );
  EDFD1 \Mem_reg[16][26]  ( .D(n24775), .E(n6471), .CP(clk), .QN(n3008) );
  EDFD1 \Mem_reg[15][26]  ( .D(n24775), .E(n6472), .CP(clk), .QN(n2960) );
  EDFD1 \Mem_reg[14][26]  ( .D(n24775), .E(n24720), .CP(clk), .QN(n2912) );
  EDFD1 \Mem_reg[13][26]  ( .D(n24775), .E(n24709), .CP(clk), .QN(n2864) );
  EDFD1 \Mem_reg[12][26]  ( .D(n24775), .E(n24717), .CP(clk), .QN(n2816) );
  EDFD1 \Mem_reg[11][26]  ( .D(n24775), .E(n24707), .CP(clk), .QN(n2768) );
  EDFD1 \Mem_reg[10][26]  ( .D(n24775), .E(n6477), .CP(clk), .QN(n2720) );
  EDFD1 \Mem_reg[9][26]  ( .D(n24775), .E(n24708), .CP(clk), .QN(n2672) );
  EDFD1 \Mem_reg[8][26]  ( .D(n24775), .E(n15642), .CP(clk), .QN(n2624) );
  EDFD1 \Mem_reg[7][26]  ( .D(n24775), .E(n24718), .CP(clk), .QN(n2576) );
  EDFD1 \Mem_reg[6][26]  ( .D(n24775), .E(n24716), .CP(clk), .QN(n2528) );
  EDFD1 \Mem_reg[5][26]  ( .D(n24775), .E(n24719), .CP(clk), .QN(n2480) );
  EDFD1 \Mem_reg[4][26]  ( .D(n24775), .E(n24706), .CP(clk), .QN(n2432) );
  EDFD1 \Mem_reg[3][26]  ( .D(n24775), .E(n24721), .CP(clk), .QN(n2384) );
  EDFD1 \Mem_reg[2][26]  ( .D(n24775), .E(n6460), .CP(clk), .QN(n2336) );
  EDFD1 \Mem_reg[1][26]  ( .D(n24775), .E(n24703), .CP(clk), .QN(n2288) );
  EDFD1 \Mem_reg[0][26]  ( .D(n24775), .E(n24705), .CP(clk), .QN(n2240) );
  EDFD1 \Mem_reg[88][25]  ( .D(n24773), .E(n6419), .CP(clk), .Q(n27137) );
  EDFD1 \Mem_reg[87][25]  ( .D(n24773), .E(n6418), .CP(clk), .QN(n6321) );
  EDFD1 \Mem_reg[86][25]  ( .D(n24773), .E(n6417), .CP(clk), .QN(n24634) );
  EDFD1 \Mem_reg[85][25]  ( .D(n24773), .E(n6416), .CP(clk), .QN(n6225) );
  EDFD1 \Mem_reg[84][25]  ( .D(n24773), .E(n6415), .CP(clk), .QN(n6177) );
  EDFD1 \Mem_reg[83][25]  ( .D(n24773), .E(n6414), .CP(clk), .QN(n6129) );
  EDFD1 \Mem_reg[82][25]  ( .D(n24773), .E(n6413), .CP(clk), .QN(n6081) );
  EDFD1 \Mem_reg[81][25]  ( .D(n24773), .E(n6412), .CP(clk), .QN(n6033) );
  EDFD1 \Mem_reg[80][25]  ( .D(n24773), .E(n6411), .CP(clk), .QN(n5985) );
  EDFD1 \Mem_reg[79][25]  ( .D(n24773), .E(n6410), .CP(clk), .QN(n5937) );
  EDFD1 \Mem_reg[78][25]  ( .D(n24773), .E(n6409), .CP(clk), .QN(n5889) );
  EDFD1 \Mem_reg[77][25]  ( .D(n24773), .E(n6408), .CP(clk), .QN(n5841) );
  EDFD1 \Mem_reg[76][25]  ( .D(n24773), .E(n6407), .CP(clk), .QN(n5793) );
  EDFD1 \Mem_reg[75][25]  ( .D(n24773), .E(n6406), .CP(clk), .QN(n27138) );
  EDFD1 \Mem_reg[74][25]  ( .D(n24773), .E(n6405), .CP(clk), .QN(n5697) );
  EDFD1 \Mem_reg[73][25]  ( .D(n24773), .E(n6404), .CP(clk), .QN(n27139) );
  EDFD1 \Mem_reg[72][25]  ( .D(n24773), .E(n6403), .CP(clk), .QN(n5601) );
  EDFD1 \Mem_reg[71][25]  ( .D(n24773), .E(n6402), .CP(clk), .QN(n5553) );
  EDFD1 \Mem_reg[70][25]  ( .D(n24773), .E(n6401), .CP(clk), .QN(n5505) );
  EDFD1 \Mem_reg[69][25]  ( .D(n24773), .E(n6400), .CP(clk), .QN(n5457) );
  EDFD1 \Mem_reg[68][25]  ( .D(n24773), .E(n6399), .CP(clk), .QN(n5409) );
  EDFD1 \Mem_reg[67][25]  ( .D(n24773), .E(n6398), .CP(clk), .QN(n5361) );
  EDFD1 \Mem_reg[66][25]  ( .D(n24773), .E(n6397), .CP(clk), .QN(n5313) );
  EDFD1 \Mem_reg[65][25]  ( .D(n24773), .E(n6396), .CP(clk), .QN(n15549) );
  EDFD1 \Mem_reg[64][25]  ( .D(n24773), .E(n6395), .CP(clk), .QN(n5217) );
  EDFD1 \Mem_reg[63][25]  ( .D(n24773), .E(n6456), .CP(clk), .QN(n5169) );
  EDFD1 \Mem_reg[62][25]  ( .D(n24773), .E(n6455), .CP(clk), .QN(n5121) );
  EDFD1 \Mem_reg[61][25]  ( .D(n24773), .E(n6454), .CP(clk), .QN(n18002) );
  EDFD1 \Mem_reg[60][25]  ( .D(n24773), .E(n6453), .CP(clk), .QN(n18001) );
  EDFD1 \Mem_reg[59][25]  ( .D(n24773), .E(n6452), .CP(clk), .QN(n4977) );
  EDFD1 \Mem_reg[58][25]  ( .D(n24773), .E(n6451), .CP(clk), .QN(n4929) );
  EDFD1 \Mem_reg[57][25]  ( .D(n24773), .E(n6450), .CP(clk), .QN(n4881) );
  EDFD1 \Mem_reg[56][25]  ( .D(n24773), .E(n6449), .CP(clk), .QN(n4833) );
  EDFD1 \Mem_reg[55][25]  ( .D(n24773), .E(n6448), .CP(clk), .QN(n4785) );
  EDFD1 \Mem_reg[54][25]  ( .D(n24773), .E(n6447), .CP(clk), .QN(n15548) );
  EDFD1 \Mem_reg[53][25]  ( .D(n24773), .E(n6446), .CP(clk), .QN(n4689) );
  EDFD1 \Mem_reg[52][25]  ( .D(n24773), .E(n6445), .CP(clk), .Q(n27136) );
  EDFD1 \Mem_reg[51][25]  ( .D(n24773), .E(n6444), .CP(clk), .QN(n4593) );
  EDFD1 \Mem_reg[50][25]  ( .D(n24773), .E(n6443), .CP(clk), .QN(n4545) );
  EDFD1 \Mem_reg[49][25]  ( .D(n24773), .E(n6442), .CP(clk), .QN(n4497) );
  EDFD1 \Mem_reg[48][25]  ( .D(n24773), .E(n6441), .CP(clk), .QN(n4449) );
  EDFD1 \Mem_reg[47][25]  ( .D(n24773), .E(n6440), .CP(clk), .QN(n4401) );
  EDFD1 \Mem_reg[46][25]  ( .D(n24773), .E(n6439), .CP(clk), .QN(n4353) );
  EDFD1 \Mem_reg[43][25]  ( .D(n24773), .E(n6438), .CP(clk), .QN(n4305) );
  EDFD1 \Mem_reg[42][25]  ( .D(n24773), .E(n6437), .CP(clk), .QN(n4257) );
  EDFD1 \Mem_reg[41][25]  ( .D(n24773), .E(n6436), .CP(clk), .QN(n4209) );
  EDFD1 \Mem_reg[40][25]  ( .D(n24773), .E(n6435), .CP(clk), .QN(n4161) );
  EDFD1 \Mem_reg[39][25]  ( .D(n24773), .E(n6434), .CP(clk), .QN(n4113) );
  EDFD1 \Mem_reg[38][25]  ( .D(n24773), .E(n6433), .CP(clk), .QN(n4065) );
  EDFD1 \Mem_reg[37][25]  ( .D(n24773), .E(n6432), .CP(clk), .QN(n4017) );
  EDFD1 \Mem_reg[36][25]  ( .D(n24773), .E(n6431), .CP(clk), .QN(n3969) );
  EDFD1 \Mem_reg[35][25]  ( .D(n24773), .E(n6430), .CP(clk), .QN(n3921) );
  EDFD1 \Mem_reg[34][25]  ( .D(n24773), .E(n6429), .CP(clk), .QN(n3873) );
  EDFD1 \Mem_reg[33][25]  ( .D(n24773), .E(n6428), .CP(clk), .QN(n3825) );
  EDFD1 \Mem_reg[32][25]  ( .D(n24773), .E(n6427), .CP(clk), .QN(n3777) );
  EDFD1 \Mem_reg[31][25]  ( .D(n24773), .E(n6426), .CP(clk), .QN(n3729) );
  EDFD1 \Mem_reg[30][25]  ( .D(n24773), .E(n6425), .CP(clk), .QN(n3681) );
  EDFD1 \Mem_reg[29][25]  ( .D(n24773), .E(n6424), .CP(clk), .QN(n3633) );
  EDFD1 \Mem_reg[28][25]  ( .D(n24773), .E(n6423), .CP(clk), .QN(n3585) );
  EDFD1 \Mem_reg[27][25]  ( .D(n24773), .E(n6422), .CP(clk), .QN(n3537) );
  EDFD1 \Mem_reg[26][25]  ( .D(n24773), .E(n6421), .CP(clk), .QN(n3489) );
  EDFD1 \Mem_reg[25][25]  ( .D(n24773), .E(n6420), .CP(clk), .QN(n3441) );
  EDFD1 \Mem_reg[24][25]  ( .D(n24773), .E(n6463), .CP(clk), .QN(n3393) );
  EDFD1 \Mem_reg[23][25]  ( .D(n24773), .E(n6464), .CP(clk), .QN(n3345) );
  EDFD1 \Mem_reg[22][25]  ( .D(n24773), .E(n6465), .CP(clk), .QN(n3297) );
  EDFD1 \Mem_reg[21][25]  ( .D(n24773), .E(n6466), .CP(clk), .QN(n3249) );
  EDFD1 \Mem_reg[20][25]  ( .D(n24773), .E(n6467), .CP(clk), .QN(n3201) );
  EDFD1 \Mem_reg[19][25]  ( .D(n24773), .E(n6468), .CP(clk), .QN(n3153) );
  EDFD1 \Mem_reg[18][25]  ( .D(n24773), .E(n6469), .CP(clk), .QN(n3105) );
  EDFD1 \Mem_reg[17][25]  ( .D(n24773), .E(n6470), .CP(clk), .QN(n3057) );
  EDFD1 \Mem_reg[16][25]  ( .D(n24773), .E(n6471), .CP(clk), .QN(n3009) );
  EDFD1 \Mem_reg[15][25]  ( .D(n24773), .E(n6472), .CP(clk), .QN(n2961) );
  EDFD1 \Mem_reg[14][25]  ( .D(n24773), .E(n24720), .CP(clk), .QN(n2913) );
  EDFD1 \Mem_reg[13][25]  ( .D(n24773), .E(n24709), .CP(clk), .QN(n2865) );
  EDFD1 \Mem_reg[12][25]  ( .D(n24773), .E(n24717), .CP(clk), .QN(n2817) );
  EDFD1 \Mem_reg[11][25]  ( .D(n24773), .E(n24707), .CP(clk), .QN(n2769) );
  EDFD1 \Mem_reg[10][25]  ( .D(n24773), .E(n6477), .CP(clk), .QN(n2721) );
  EDFD1 \Mem_reg[9][25]  ( .D(n24773), .E(n24708), .CP(clk), .QN(n2673) );
  EDFD1 \Mem_reg[8][25]  ( .D(n24773), .E(n15642), .CP(clk), .QN(n2625) );
  EDFD1 \Mem_reg[7][25]  ( .D(n24773), .E(n24718), .CP(clk), .QN(n2577) );
  EDFD1 \Mem_reg[6][25]  ( .D(n24773), .E(n24716), .CP(clk), .QN(n2529) );
  EDFD1 \Mem_reg[5][25]  ( .D(n24773), .E(n24719), .CP(clk), .QN(n2481) );
  EDFD1 \Mem_reg[4][25]  ( .D(n24773), .E(n24706), .CP(clk), .QN(n2433) );
  EDFD1 \Mem_reg[3][25]  ( .D(n24773), .E(n24721), .CP(clk), .QN(n2385) );
  EDFD1 \Mem_reg[2][25]  ( .D(n24773), .E(n6460), .CP(clk), .QN(n2337) );
  EDFD1 \Mem_reg[1][25]  ( .D(n24773), .E(n24703), .CP(clk), .QN(n2289) );
  EDFD1 \Mem_reg[0][25]  ( .D(n24773), .E(n24705), .CP(clk), .QN(n2241) );
  EDFD1 \Mem_reg[88][24]  ( .D(n24771), .E(n6419), .CP(clk), .Q(n27133) );
  EDFD1 \Mem_reg[87][24]  ( .D(n24771), .E(n6418), .CP(clk), .QN(n6322) );
  EDFD1 \Mem_reg[86][24]  ( .D(n24771), .E(n6417), .CP(clk), .QN(n24631) );
  EDFD1 \Mem_reg[85][24]  ( .D(n24771), .E(n6416), .CP(clk), .QN(n6226) );
  EDFD1 \Mem_reg[84][24]  ( .D(n24771), .E(n6415), .CP(clk), .QN(n6178) );
  EDFD1 \Mem_reg[83][24]  ( .D(n24771), .E(n6414), .CP(clk), .QN(n6130) );
  EDFD1 \Mem_reg[82][24]  ( .D(n24771), .E(n6413), .CP(clk), .QN(n6082) );
  EDFD1 \Mem_reg[81][24]  ( .D(n24771), .E(n6412), .CP(clk), .QN(n6034) );
  EDFD1 \Mem_reg[80][24]  ( .D(n24771), .E(n6411), .CP(clk), .QN(n5986) );
  EDFD1 \Mem_reg[79][24]  ( .D(n24771), .E(n6410), .CP(clk), .QN(n5938) );
  EDFD1 \Mem_reg[78][24]  ( .D(n24771), .E(n6409), .CP(clk), .QN(n5890) );
  EDFD1 \Mem_reg[77][24]  ( .D(n24771), .E(n6408), .CP(clk), .QN(n5842) );
  EDFD1 \Mem_reg[76][24]  ( .D(n24771), .E(n6407), .CP(clk), .QN(n5794) );
  EDFD1 \Mem_reg[75][24]  ( .D(n24771), .E(n6406), .CP(clk), .QN(n27134) );
  EDFD1 \Mem_reg[74][24]  ( .D(n24771), .E(n6405), .CP(clk), .QN(n5698) );
  EDFD1 \Mem_reg[73][24]  ( .D(n24771), .E(n6404), .CP(clk), .QN(n27135) );
  EDFD1 \Mem_reg[72][24]  ( .D(n24771), .E(n6403), .CP(clk), .QN(n5602) );
  EDFD1 \Mem_reg[71][24]  ( .D(n24771), .E(n6402), .CP(clk), .QN(n5554) );
  EDFD1 \Mem_reg[70][24]  ( .D(n24771), .E(n6401), .CP(clk), .QN(n5506) );
  EDFD1 \Mem_reg[69][24]  ( .D(n24771), .E(n6400), .CP(clk), .QN(n5458) );
  EDFD1 \Mem_reg[68][24]  ( .D(n24771), .E(n6399), .CP(clk), .QN(n5410) );
  EDFD1 \Mem_reg[67][24]  ( .D(n24771), .E(n6398), .CP(clk), .QN(n5362) );
  EDFD1 \Mem_reg[66][24]  ( .D(n24771), .E(n6397), .CP(clk), .QN(n5314) );
  EDFD1 \Mem_reg[65][24]  ( .D(n24771), .E(n6396), .CP(clk), .QN(n15545) );
  EDFD1 \Mem_reg[64][24]  ( .D(n24771), .E(n6395), .CP(clk), .QN(n5218) );
  EDFD1 \Mem_reg[63][24]  ( .D(n24771), .E(n6456), .CP(clk), .QN(n5170) );
  EDFD1 \Mem_reg[62][24]  ( .D(n24771), .E(n6455), .CP(clk), .QN(n5122) );
  EDFD1 \Mem_reg[61][24]  ( .D(n24771), .E(n6454), .CP(clk), .QN(n17999) );
  EDFD1 \Mem_reg[60][24]  ( .D(n24771), .E(n6453), .CP(clk), .QN(n17998) );
  EDFD1 \Mem_reg[59][24]  ( .D(n24771), .E(n6452), .CP(clk), .QN(n4978) );
  EDFD1 \Mem_reg[58][24]  ( .D(n24771), .E(n6451), .CP(clk), .QN(n4930) );
  EDFD1 \Mem_reg[57][24]  ( .D(n24771), .E(n6450), .CP(clk), .QN(n4882) );
  EDFD1 \Mem_reg[56][24]  ( .D(n24771), .E(n6449), .CP(clk), .QN(n4834) );
  EDFD1 \Mem_reg[55][24]  ( .D(n24771), .E(n6448), .CP(clk), .QN(n4786) );
  EDFD1 \Mem_reg[54][24]  ( .D(n24771), .E(n6447), .CP(clk), .QN(n15544) );
  EDFD1 \Mem_reg[53][24]  ( .D(n24771), .E(n6446), .CP(clk), .QN(n4690) );
  EDFD1 \Mem_reg[52][24]  ( .D(n24771), .E(n6445), .CP(clk), .Q(n27132) );
  EDFD1 \Mem_reg[51][24]  ( .D(n24771), .E(n6444), .CP(clk), .QN(n4594) );
  EDFD1 \Mem_reg[50][24]  ( .D(n24771), .E(n6443), .CP(clk), .QN(n4546) );
  EDFD1 \Mem_reg[49][24]  ( .D(n24771), .E(n6442), .CP(clk), .QN(n4498) );
  EDFD1 \Mem_reg[48][24]  ( .D(n24771), .E(n6441), .CP(clk), .QN(n4450) );
  EDFD1 \Mem_reg[47][24]  ( .D(n24771), .E(n6440), .CP(clk), .QN(n4402) );
  EDFD1 \Mem_reg[46][24]  ( .D(n24771), .E(n6439), .CP(clk), .QN(n4354) );
  EDFD1 \Mem_reg[43][24]  ( .D(n24771), .E(n6438), .CP(clk), .QN(n4306) );
  EDFD1 \Mem_reg[42][24]  ( .D(n24771), .E(n6437), .CP(clk), .QN(n4258) );
  EDFD1 \Mem_reg[41][24]  ( .D(n24771), .E(n6436), .CP(clk), .QN(n4210) );
  EDFD1 \Mem_reg[40][24]  ( .D(n24771), .E(n6435), .CP(clk), .QN(n4162) );
  EDFD1 \Mem_reg[39][24]  ( .D(n24771), .E(n6434), .CP(clk), .QN(n4114) );
  EDFD1 \Mem_reg[38][24]  ( .D(n24771), .E(n6433), .CP(clk), .QN(n4066) );
  EDFD1 \Mem_reg[37][24]  ( .D(n24771), .E(n6432), .CP(clk), .QN(n4018) );
  EDFD1 \Mem_reg[36][24]  ( .D(n24771), .E(n6431), .CP(clk), .QN(n3970) );
  EDFD1 \Mem_reg[35][24]  ( .D(n24771), .E(n6430), .CP(clk), .QN(n3922) );
  EDFD1 \Mem_reg[34][24]  ( .D(n24771), .E(n6429), .CP(clk), .QN(n3874) );
  EDFD1 \Mem_reg[33][24]  ( .D(n24771), .E(n6428), .CP(clk), .QN(n3826) );
  EDFD1 \Mem_reg[32][24]  ( .D(n24771), .E(n6427), .CP(clk), .QN(n3778) );
  EDFD1 \Mem_reg[31][24]  ( .D(n24771), .E(n6426), .CP(clk), .QN(n3730) );
  EDFD1 \Mem_reg[30][24]  ( .D(n24771), .E(n6425), .CP(clk), .QN(n3682) );
  EDFD1 \Mem_reg[29][24]  ( .D(n24771), .E(n6424), .CP(clk), .QN(n3634) );
  EDFD1 \Mem_reg[28][24]  ( .D(n24771), .E(n6423), .CP(clk), .QN(n3586) );
  EDFD1 \Mem_reg[27][24]  ( .D(n24771), .E(n6422), .CP(clk), .QN(n3538) );
  EDFD1 \Mem_reg[26][24]  ( .D(n24771), .E(n6421), .CP(clk), .QN(n3490) );
  EDFD1 \Mem_reg[25][24]  ( .D(n24771), .E(n6420), .CP(clk), .QN(n3442) );
  EDFD1 \Mem_reg[24][24]  ( .D(n24771), .E(n6463), .CP(clk), .QN(n3394) );
  EDFD1 \Mem_reg[23][24]  ( .D(n24771), .E(n6464), .CP(clk), .QN(n3346) );
  EDFD1 \Mem_reg[22][24]  ( .D(n24771), .E(n6465), .CP(clk), .QN(n3298) );
  EDFD1 \Mem_reg[21][24]  ( .D(n24771), .E(n6466), .CP(clk), .QN(n3250) );
  EDFD1 \Mem_reg[20][24]  ( .D(n24771), .E(n6467), .CP(clk), .QN(n3202) );
  EDFD1 \Mem_reg[19][24]  ( .D(n24771), .E(n6468), .CP(clk), .QN(n3154) );
  EDFD1 \Mem_reg[18][24]  ( .D(n24771), .E(n6469), .CP(clk), .QN(n3106) );
  EDFD1 \Mem_reg[17][24]  ( .D(n24771), .E(n6470), .CP(clk), .QN(n3058) );
  EDFD1 \Mem_reg[16][24]  ( .D(n24771), .E(n6471), .CP(clk), .QN(n3010) );
  EDFD1 \Mem_reg[15][24]  ( .D(n24771), .E(n6472), .CP(clk), .QN(n2962) );
  EDFD1 \Mem_reg[14][24]  ( .D(n24771), .E(n24720), .CP(clk), .QN(n2914) );
  EDFD1 \Mem_reg[13][24]  ( .D(n24771), .E(n24709), .CP(clk), .QN(n2866) );
  EDFD1 \Mem_reg[12][24]  ( .D(n24771), .E(n24717), .CP(clk), .QN(n2818) );
  EDFD1 \Mem_reg[11][24]  ( .D(n24771), .E(n24707), .CP(clk), .QN(n2770) );
  EDFD1 \Mem_reg[10][24]  ( .D(n24771), .E(n6477), .CP(clk), .QN(n2722) );
  EDFD1 \Mem_reg[9][24]  ( .D(n24771), .E(n24708), .CP(clk), .QN(n2674) );
  EDFD1 \Mem_reg[8][24]  ( .D(n24771), .E(n15642), .CP(clk), .QN(n2626) );
  EDFD1 \Mem_reg[7][24]  ( .D(n24771), .E(n24718), .CP(clk), .QN(n2578) );
  EDFD1 \Mem_reg[6][24]  ( .D(n24771), .E(n24716), .CP(clk), .QN(n2530) );
  EDFD1 \Mem_reg[5][24]  ( .D(n24771), .E(n24719), .CP(clk), .QN(n2482) );
  EDFD1 \Mem_reg[4][24]  ( .D(n24771), .E(n24706), .CP(clk), .QN(n2434) );
  EDFD1 \Mem_reg[3][24]  ( .D(n24771), .E(n24721), .CP(clk), .QN(n2386) );
  EDFD1 \Mem_reg[2][24]  ( .D(n24771), .E(n6460), .CP(clk), .QN(n2338) );
  EDFD1 \Mem_reg[1][24]  ( .D(n24771), .E(n24703), .CP(clk), .QN(n2290) );
  EDFD1 \Mem_reg[0][24]  ( .D(n24771), .E(n24705), .CP(clk), .QN(n2242) );
  EDFD1 \Mem_reg[88][23]  ( .D(n24769), .E(n6419), .CP(clk), .Q(n27129) );
  EDFD1 \Mem_reg[87][23]  ( .D(n24769), .E(n6418), .CP(clk), .QN(n6323) );
  EDFD1 \Mem_reg[86][23]  ( .D(n24769), .E(n6417), .CP(clk), .QN(n24628) );
  EDFD1 \Mem_reg[85][23]  ( .D(n24769), .E(n6416), .CP(clk), .QN(n6227) );
  EDFD1 \Mem_reg[84][23]  ( .D(n24769), .E(n6415), .CP(clk), .QN(n6179) );
  EDFD1 \Mem_reg[83][23]  ( .D(n24769), .E(n6414), .CP(clk), .QN(n6131) );
  EDFD1 \Mem_reg[82][23]  ( .D(n24769), .E(n6413), .CP(clk), .QN(n6083) );
  EDFD1 \Mem_reg[81][23]  ( .D(n24769), .E(n6412), .CP(clk), .QN(n6035) );
  EDFD1 \Mem_reg[80][23]  ( .D(n24769), .E(n6411), .CP(clk), .QN(n5987) );
  EDFD1 \Mem_reg[79][23]  ( .D(n24769), .E(n6410), .CP(clk), .QN(n5939) );
  EDFD1 \Mem_reg[78][23]  ( .D(n24769), .E(n6409), .CP(clk), .QN(n5891) );
  EDFD1 \Mem_reg[77][23]  ( .D(n24769), .E(n6408), .CP(clk), .QN(n5843) );
  EDFD1 \Mem_reg[76][23]  ( .D(n24769), .E(n6407), .CP(clk), .QN(n5795) );
  EDFD1 \Mem_reg[75][23]  ( .D(n24769), .E(n6406), .CP(clk), .QN(n27130) );
  EDFD1 \Mem_reg[74][23]  ( .D(n24769), .E(n6405), .CP(clk), .QN(n5699) );
  EDFD1 \Mem_reg[73][23]  ( .D(n24769), .E(n6404), .CP(clk), .QN(n27131) );
  EDFD1 \Mem_reg[72][23]  ( .D(n24769), .E(n6403), .CP(clk), .QN(n5603) );
  EDFD1 \Mem_reg[71][23]  ( .D(n24769), .E(n6402), .CP(clk), .QN(n5555) );
  EDFD1 \Mem_reg[70][23]  ( .D(n24769), .E(n6401), .CP(clk), .QN(n5507) );
  EDFD1 \Mem_reg[69][23]  ( .D(n24769), .E(n6400), .CP(clk), .QN(n5459) );
  EDFD1 \Mem_reg[68][23]  ( .D(n24769), .E(n6399), .CP(clk), .QN(n5411) );
  EDFD1 \Mem_reg[67][23]  ( .D(n24769), .E(n6398), .CP(clk), .QN(n5363) );
  EDFD1 \Mem_reg[66][23]  ( .D(n24769), .E(n6397), .CP(clk), .QN(n5315) );
  EDFD1 \Mem_reg[65][23]  ( .D(n24769), .E(n6396), .CP(clk), .QN(n15541) );
  EDFD1 \Mem_reg[64][23]  ( .D(n24769), .E(n6395), .CP(clk), .QN(n5219) );
  EDFD1 \Mem_reg[63][23]  ( .D(n24769), .E(n6456), .CP(clk), .QN(n5171) );
  EDFD1 \Mem_reg[62][23]  ( .D(n24769), .E(n6455), .CP(clk), .QN(n5123) );
  EDFD1 \Mem_reg[61][23]  ( .D(n24769), .E(n6454), .CP(clk), .QN(n17996) );
  EDFD1 \Mem_reg[60][23]  ( .D(n24769), .E(n6453), .CP(clk), .QN(n17995) );
  EDFD1 \Mem_reg[59][23]  ( .D(n24769), .E(n6452), .CP(clk), .QN(n4979) );
  EDFD1 \Mem_reg[58][23]  ( .D(n24769), .E(n6451), .CP(clk), .QN(n4931) );
  EDFD1 \Mem_reg[57][23]  ( .D(n24769), .E(n6450), .CP(clk), .QN(n4883) );
  EDFD1 \Mem_reg[56][23]  ( .D(n24769), .E(n6449), .CP(clk), .QN(n4835) );
  EDFD1 \Mem_reg[55][23]  ( .D(n24769), .E(n6448), .CP(clk), .QN(n4787) );
  EDFD1 \Mem_reg[54][23]  ( .D(n24769), .E(n6447), .CP(clk), .QN(n15540) );
  EDFD1 \Mem_reg[53][23]  ( .D(n24769), .E(n6446), .CP(clk), .QN(n4691) );
  EDFD1 \Mem_reg[52][23]  ( .D(n24769), .E(n6445), .CP(clk), .Q(n27128) );
  EDFD1 \Mem_reg[51][23]  ( .D(n24769), .E(n6444), .CP(clk), .QN(n4595) );
  EDFD1 \Mem_reg[50][23]  ( .D(n24769), .E(n6443), .CP(clk), .QN(n4547) );
  EDFD1 \Mem_reg[49][23]  ( .D(n24769), .E(n6442), .CP(clk), .QN(n4499) );
  EDFD1 \Mem_reg[48][23]  ( .D(n24769), .E(n6441), .CP(clk), .QN(n4451) );
  EDFD1 \Mem_reg[47][23]  ( .D(n24769), .E(n6440), .CP(clk), .QN(n4403) );
  EDFD1 \Mem_reg[46][23]  ( .D(n24769), .E(n6439), .CP(clk), .QN(n4355) );
  EDFD1 \Mem_reg[43][23]  ( .D(n24769), .E(n6438), .CP(clk), .QN(n4307) );
  EDFD1 \Mem_reg[42][23]  ( .D(n24769), .E(n6437), .CP(clk), .QN(n4259) );
  EDFD1 \Mem_reg[41][23]  ( .D(n24769), .E(n6436), .CP(clk), .QN(n4211) );
  EDFD1 \Mem_reg[40][23]  ( .D(n24769), .E(n6435), .CP(clk), .QN(n4163) );
  EDFD1 \Mem_reg[39][23]  ( .D(n24769), .E(n6434), .CP(clk), .QN(n4115) );
  EDFD1 \Mem_reg[38][23]  ( .D(n24769), .E(n6433), .CP(clk), .QN(n4067) );
  EDFD1 \Mem_reg[37][23]  ( .D(n24769), .E(n6432), .CP(clk), .QN(n4019) );
  EDFD1 \Mem_reg[36][23]  ( .D(n24769), .E(n6431), .CP(clk), .QN(n3971) );
  EDFD1 \Mem_reg[35][23]  ( .D(n24769), .E(n6430), .CP(clk), .QN(n3923) );
  EDFD1 \Mem_reg[34][23]  ( .D(n24769), .E(n6429), .CP(clk), .QN(n3875) );
  EDFD1 \Mem_reg[33][23]  ( .D(n24769), .E(n6428), .CP(clk), .QN(n3827) );
  EDFD1 \Mem_reg[32][23]  ( .D(n24769), .E(n6427), .CP(clk), .QN(n3779) );
  EDFD1 \Mem_reg[31][23]  ( .D(n24769), .E(n6426), .CP(clk), .QN(n3731) );
  EDFD1 \Mem_reg[30][23]  ( .D(n24769), .E(n6425), .CP(clk), .QN(n3683) );
  EDFD1 \Mem_reg[29][23]  ( .D(n24769), .E(n6424), .CP(clk), .QN(n3635) );
  EDFD1 \Mem_reg[28][23]  ( .D(n24769), .E(n6423), .CP(clk), .QN(n3587) );
  EDFD1 \Mem_reg[27][23]  ( .D(n24769), .E(n6422), .CP(clk), .QN(n3539) );
  EDFD1 \Mem_reg[26][23]  ( .D(n24769), .E(n6421), .CP(clk), .QN(n3491) );
  EDFD1 \Mem_reg[25][23]  ( .D(n24769), .E(n6420), .CP(clk), .QN(n3443) );
  EDFD1 \Mem_reg[24][23]  ( .D(n24769), .E(n6463), .CP(clk), .QN(n3395) );
  EDFD1 \Mem_reg[23][23]  ( .D(n24769), .E(n6464), .CP(clk), .QN(n3347) );
  EDFD1 \Mem_reg[22][23]  ( .D(n24769), .E(n6465), .CP(clk), .QN(n3299) );
  EDFD1 \Mem_reg[21][23]  ( .D(n24769), .E(n6466), .CP(clk), .QN(n3251) );
  EDFD1 \Mem_reg[20][23]  ( .D(n24769), .E(n6467), .CP(clk), .QN(n3203) );
  EDFD1 \Mem_reg[19][23]  ( .D(n24769), .E(n6468), .CP(clk), .QN(n3155) );
  EDFD1 \Mem_reg[18][23]  ( .D(n24769), .E(n6469), .CP(clk), .QN(n3107) );
  EDFD1 \Mem_reg[17][23]  ( .D(n24769), .E(n6470), .CP(clk), .QN(n3059) );
  EDFD1 \Mem_reg[16][23]  ( .D(n24769), .E(n6471), .CP(clk), .QN(n3011) );
  EDFD1 \Mem_reg[15][23]  ( .D(n24769), .E(n6472), .CP(clk), .QN(n2963) );
  EDFD1 \Mem_reg[14][23]  ( .D(n24769), .E(n24720), .CP(clk), .QN(n2915) );
  EDFD1 \Mem_reg[13][23]  ( .D(n24769), .E(n24709), .CP(clk), .QN(n2867) );
  EDFD1 \Mem_reg[12][23]  ( .D(n24769), .E(n24717), .CP(clk), .QN(n2819) );
  EDFD1 \Mem_reg[11][23]  ( .D(n24769), .E(n24707), .CP(clk), .QN(n2771) );
  EDFD1 \Mem_reg[10][23]  ( .D(n24769), .E(n6477), .CP(clk), .QN(n2723) );
  EDFD1 \Mem_reg[9][23]  ( .D(n24769), .E(n24708), .CP(clk), .QN(n2675) );
  EDFD1 \Mem_reg[8][23]  ( .D(n24769), .E(n15642), .CP(clk), .QN(n2627) );
  EDFD1 \Mem_reg[7][23]  ( .D(n24769), .E(n24718), .CP(clk), .QN(n2579) );
  EDFD1 \Mem_reg[6][23]  ( .D(n24769), .E(n24716), .CP(clk), .QN(n2531) );
  EDFD1 \Mem_reg[5][23]  ( .D(n24769), .E(n24719), .CP(clk), .QN(n2483) );
  EDFD1 \Mem_reg[4][23]  ( .D(n24769), .E(n24706), .CP(clk), .QN(n2435) );
  EDFD1 \Mem_reg[3][23]  ( .D(n24769), .E(n24721), .CP(clk), .QN(n2387) );
  EDFD1 \Mem_reg[2][23]  ( .D(n24769), .E(n6460), .CP(clk), .QN(n2339) );
  EDFD1 \Mem_reg[1][23]  ( .D(n24769), .E(n24703), .CP(clk), .QN(n2291) );
  EDFD1 \Mem_reg[0][23]  ( .D(n24769), .E(n24705), .CP(clk), .QN(n2243) );
  EDFD1 \Mem_reg[88][22]  ( .D(n24767), .E(n6419), .CP(clk), .Q(n27125) );
  EDFD1 \Mem_reg[87][22]  ( .D(n24767), .E(n6418), .CP(clk), .QN(n6324) );
  EDFD1 \Mem_reg[86][22]  ( .D(n24767), .E(n6417), .CP(clk), .QN(n24625) );
  EDFD1 \Mem_reg[85][22]  ( .D(n24767), .E(n6416), .CP(clk), .QN(n6228) );
  EDFD1 \Mem_reg[84][22]  ( .D(n24767), .E(n6415), .CP(clk), .QN(n6180) );
  EDFD1 \Mem_reg[83][22]  ( .D(n24767), .E(n6414), .CP(clk), .QN(n6132) );
  EDFD1 \Mem_reg[82][22]  ( .D(n24767), .E(n6413), .CP(clk), .QN(n6084) );
  EDFD1 \Mem_reg[81][22]  ( .D(n24767), .E(n6412), .CP(clk), .QN(n6036) );
  EDFD1 \Mem_reg[80][22]  ( .D(n24767), .E(n6411), .CP(clk), .QN(n5988) );
  EDFD1 \Mem_reg[79][22]  ( .D(n24767), .E(n6410), .CP(clk), .QN(n5940) );
  EDFD1 \Mem_reg[78][22]  ( .D(n24767), .E(n6409), .CP(clk), .QN(n5892) );
  EDFD1 \Mem_reg[77][22]  ( .D(n24767), .E(n6408), .CP(clk), .QN(n5844) );
  EDFD1 \Mem_reg[76][22]  ( .D(n24767), .E(n6407), .CP(clk), .QN(n5796) );
  EDFD1 \Mem_reg[75][22]  ( .D(n24767), .E(n6406), .CP(clk), .QN(n27126) );
  EDFD1 \Mem_reg[74][22]  ( .D(n24767), .E(n6405), .CP(clk), .QN(n5700) );
  EDFD1 \Mem_reg[73][22]  ( .D(n24767), .E(n6404), .CP(clk), .QN(n27127) );
  EDFD1 \Mem_reg[72][22]  ( .D(n24767), .E(n6403), .CP(clk), .QN(n5604) );
  EDFD1 \Mem_reg[71][22]  ( .D(n24767), .E(n6402), .CP(clk), .QN(n5556) );
  EDFD1 \Mem_reg[70][22]  ( .D(n24767), .E(n6401), .CP(clk), .QN(n5508) );
  EDFD1 \Mem_reg[69][22]  ( .D(n24767), .E(n6400), .CP(clk), .QN(n5460) );
  EDFD1 \Mem_reg[68][22]  ( .D(n24767), .E(n6399), .CP(clk), .QN(n5412) );
  EDFD1 \Mem_reg[67][22]  ( .D(n24767), .E(n6398), .CP(clk), .QN(n5364) );
  EDFD1 \Mem_reg[66][22]  ( .D(n24767), .E(n6397), .CP(clk), .QN(n5316) );
  EDFD1 \Mem_reg[65][22]  ( .D(n24767), .E(n6396), .CP(clk), .QN(n15537) );
  EDFD1 \Mem_reg[64][22]  ( .D(n24767), .E(n6395), .CP(clk), .QN(n5220) );
  EDFD1 \Mem_reg[63][22]  ( .D(n24767), .E(n6456), .CP(clk), .QN(n5172) );
  EDFD1 \Mem_reg[62][22]  ( .D(n24767), .E(n6455), .CP(clk), .QN(n5124) );
  EDFD1 \Mem_reg[61][22]  ( .D(n24767), .E(n6454), .CP(clk), .QN(n17993) );
  EDFD1 \Mem_reg[60][22]  ( .D(n24767), .E(n6453), .CP(clk), .QN(n17992) );
  EDFD1 \Mem_reg[59][22]  ( .D(n24767), .E(n6452), .CP(clk), .QN(n4980) );
  EDFD1 \Mem_reg[58][22]  ( .D(n24767), .E(n6451), .CP(clk), .QN(n4932) );
  EDFD1 \Mem_reg[57][22]  ( .D(n24767), .E(n6450), .CP(clk), .QN(n4884) );
  EDFD1 \Mem_reg[56][22]  ( .D(n24767), .E(n6449), .CP(clk), .QN(n4836) );
  EDFD1 \Mem_reg[55][22]  ( .D(n24767), .E(n6448), .CP(clk), .QN(n4788) );
  EDFD1 \Mem_reg[54][22]  ( .D(n24767), .E(n6447), .CP(clk), .QN(n15536) );
  EDFD1 \Mem_reg[53][22]  ( .D(n24767), .E(n6446), .CP(clk), .QN(n4692) );
  EDFD1 \Mem_reg[52][22]  ( .D(n24767), .E(n6445), .CP(clk), .Q(n27124) );
  EDFD1 \Mem_reg[51][22]  ( .D(n24767), .E(n6444), .CP(clk), .QN(n4596) );
  EDFD1 \Mem_reg[50][22]  ( .D(n24767), .E(n6443), .CP(clk), .QN(n4548) );
  EDFD1 \Mem_reg[49][22]  ( .D(n24767), .E(n6442), .CP(clk), .QN(n4500) );
  EDFD1 \Mem_reg[48][22]  ( .D(n24767), .E(n6441), .CP(clk), .QN(n4452) );
  EDFD1 \Mem_reg[47][22]  ( .D(n24767), .E(n6440), .CP(clk), .QN(n4404) );
  EDFD1 \Mem_reg[46][22]  ( .D(n24767), .E(n6439), .CP(clk), .QN(n4356) );
  EDFD1 \Mem_reg[43][22]  ( .D(n24767), .E(n6438), .CP(clk), .QN(n4308) );
  EDFD1 \Mem_reg[42][22]  ( .D(n24767), .E(n6437), .CP(clk), .QN(n4260) );
  EDFD1 \Mem_reg[41][22]  ( .D(n24767), .E(n6436), .CP(clk), .QN(n4212) );
  EDFD1 \Mem_reg[40][22]  ( .D(n24767), .E(n6435), .CP(clk), .QN(n4164) );
  EDFD1 \Mem_reg[39][22]  ( .D(n24767), .E(n6434), .CP(clk), .QN(n4116) );
  EDFD1 \Mem_reg[38][22]  ( .D(n24767), .E(n6433), .CP(clk), .QN(n4068) );
  EDFD1 \Mem_reg[37][22]  ( .D(n24767), .E(n6432), .CP(clk), .QN(n4020) );
  EDFD1 \Mem_reg[36][22]  ( .D(n24767), .E(n6431), .CP(clk), .QN(n3972) );
  EDFD1 \Mem_reg[35][22]  ( .D(n24767), .E(n6430), .CP(clk), .QN(n3924) );
  EDFD1 \Mem_reg[34][22]  ( .D(n24767), .E(n6429), .CP(clk), .QN(n3876) );
  EDFD1 \Mem_reg[33][22]  ( .D(n24767), .E(n6428), .CP(clk), .QN(n3828) );
  EDFD1 \Mem_reg[32][22]  ( .D(n24767), .E(n6427), .CP(clk), .QN(n3780) );
  EDFD1 \Mem_reg[31][22]  ( .D(n24767), .E(n6426), .CP(clk), .QN(n3732) );
  EDFD1 \Mem_reg[30][22]  ( .D(n24767), .E(n6425), .CP(clk), .QN(n3684) );
  EDFD1 \Mem_reg[29][22]  ( .D(n24767), .E(n6424), .CP(clk), .QN(n3636) );
  EDFD1 \Mem_reg[28][22]  ( .D(n24767), .E(n6423), .CP(clk), .QN(n3588) );
  EDFD1 \Mem_reg[27][22]  ( .D(n24767), .E(n6422), .CP(clk), .QN(n3540) );
  EDFD1 \Mem_reg[26][22]  ( .D(n24767), .E(n6421), .CP(clk), .QN(n3492) );
  EDFD1 \Mem_reg[25][22]  ( .D(n24767), .E(n6420), .CP(clk), .QN(n3444) );
  EDFD1 \Mem_reg[24][22]  ( .D(n24767), .E(n6463), .CP(clk), .QN(n3396) );
  EDFD1 \Mem_reg[23][22]  ( .D(n24767), .E(n6464), .CP(clk), .QN(n3348) );
  EDFD1 \Mem_reg[22][22]  ( .D(n24767), .E(n6465), .CP(clk), .QN(n3300) );
  EDFD1 \Mem_reg[21][22]  ( .D(n24767), .E(n6466), .CP(clk), .QN(n3252) );
  EDFD1 \Mem_reg[20][22]  ( .D(n24767), .E(n6467), .CP(clk), .QN(n3204) );
  EDFD1 \Mem_reg[19][22]  ( .D(n24767), .E(n6468), .CP(clk), .QN(n3156) );
  EDFD1 \Mem_reg[18][22]  ( .D(n24767), .E(n6469), .CP(clk), .QN(n3108) );
  EDFD1 \Mem_reg[17][22]  ( .D(n24767), .E(n6470), .CP(clk), .QN(n3060) );
  EDFD1 \Mem_reg[16][22]  ( .D(n24767), .E(n6471), .CP(clk), .QN(n3012) );
  EDFD1 \Mem_reg[15][22]  ( .D(n24767), .E(n6472), .CP(clk), .QN(n2964) );
  EDFD1 \Mem_reg[14][22]  ( .D(n24767), .E(n24720), .CP(clk), .QN(n2916) );
  EDFD1 \Mem_reg[13][22]  ( .D(n24767), .E(n24709), .CP(clk), .QN(n2868) );
  EDFD1 \Mem_reg[12][22]  ( .D(n24767), .E(n24717), .CP(clk), .QN(n2820) );
  EDFD1 \Mem_reg[11][22]  ( .D(n24767), .E(n24707), .CP(clk), .QN(n2772) );
  EDFD1 \Mem_reg[10][22]  ( .D(n24767), .E(n6477), .CP(clk), .QN(n2724) );
  EDFD1 \Mem_reg[9][22]  ( .D(n24767), .E(n24708), .CP(clk), .QN(n2676) );
  EDFD1 \Mem_reg[8][22]  ( .D(n24767), .E(n15642), .CP(clk), .QN(n2628) );
  EDFD1 \Mem_reg[7][22]  ( .D(n24767), .E(n24718), .CP(clk), .QN(n2580) );
  EDFD1 \Mem_reg[6][22]  ( .D(n24767), .E(n24716), .CP(clk), .QN(n2532) );
  EDFD1 \Mem_reg[5][22]  ( .D(n24767), .E(n24719), .CP(clk), .QN(n2484) );
  EDFD1 \Mem_reg[4][22]  ( .D(n24767), .E(n24706), .CP(clk), .QN(n2436) );
  EDFD1 \Mem_reg[3][22]  ( .D(n24767), .E(n24721), .CP(clk), .QN(n2388) );
  EDFD1 \Mem_reg[2][22]  ( .D(n24767), .E(n6460), .CP(clk), .QN(n2340) );
  EDFD1 \Mem_reg[1][22]  ( .D(n24767), .E(n24703), .CP(clk), .QN(n2292) );
  EDFD1 \Mem_reg[0][22]  ( .D(n24767), .E(n24705), .CP(clk), .QN(n2244) );
  EDFD1 \Mem_reg[88][21]  ( .D(n24765), .E(n6419), .CP(clk), .Q(n27121) );
  EDFD1 \Mem_reg[87][21]  ( .D(n24765), .E(n6418), .CP(clk), .QN(n6325) );
  EDFD1 \Mem_reg[86][21]  ( .D(n24765), .E(n6417), .CP(clk), .QN(n24622) );
  EDFD1 \Mem_reg[85][21]  ( .D(n24765), .E(n6416), .CP(clk), .QN(n6229) );
  EDFD1 \Mem_reg[84][21]  ( .D(n24765), .E(n6415), .CP(clk), .QN(n6181) );
  EDFD1 \Mem_reg[83][21]  ( .D(n24765), .E(n6414), .CP(clk), .QN(n6133) );
  EDFD1 \Mem_reg[82][21]  ( .D(n24765), .E(n6413), .CP(clk), .QN(n6085) );
  EDFD1 \Mem_reg[81][21]  ( .D(n24765), .E(n6412), .CP(clk), .QN(n6037) );
  EDFD1 \Mem_reg[80][21]  ( .D(n24765), .E(n6411), .CP(clk), .QN(n5989) );
  EDFD1 \Mem_reg[79][21]  ( .D(n24765), .E(n6410), .CP(clk), .QN(n5941) );
  EDFD1 \Mem_reg[78][21]  ( .D(n24765), .E(n6409), .CP(clk), .QN(n5893) );
  EDFD1 \Mem_reg[77][21]  ( .D(n24765), .E(n6408), .CP(clk), .QN(n5845) );
  EDFD1 \Mem_reg[76][21]  ( .D(n24765), .E(n6407), .CP(clk), .QN(n5797) );
  EDFD1 \Mem_reg[75][21]  ( .D(n24765), .E(n6406), .CP(clk), .QN(n27122) );
  EDFD1 \Mem_reg[74][21]  ( .D(n24765), .E(n6405), .CP(clk), .QN(n5701) );
  EDFD1 \Mem_reg[73][21]  ( .D(n24765), .E(n6404), .CP(clk), .QN(n27123) );
  EDFD1 \Mem_reg[72][21]  ( .D(n24765), .E(n6403), .CP(clk), .QN(n5605) );
  EDFD1 \Mem_reg[71][21]  ( .D(n24765), .E(n6402), .CP(clk), .QN(n5557) );
  EDFD1 \Mem_reg[70][21]  ( .D(n24765), .E(n6401), .CP(clk), .QN(n5509) );
  EDFD1 \Mem_reg[69][21]  ( .D(n24765), .E(n6400), .CP(clk), .QN(n5461) );
  EDFD1 \Mem_reg[68][21]  ( .D(n24765), .E(n6399), .CP(clk), .QN(n5413) );
  EDFD1 \Mem_reg[67][21]  ( .D(n24765), .E(n6398), .CP(clk), .QN(n5365) );
  EDFD1 \Mem_reg[66][21]  ( .D(n24765), .E(n6397), .CP(clk), .QN(n5317) );
  EDFD1 \Mem_reg[65][21]  ( .D(n24765), .E(n6396), .CP(clk), .QN(n15533) );
  EDFD1 \Mem_reg[64][21]  ( .D(n24765), .E(n6395), .CP(clk), .QN(n5221) );
  EDFD1 \Mem_reg[63][21]  ( .D(n24765), .E(n6456), .CP(clk), .QN(n5173) );
  EDFD1 \Mem_reg[62][21]  ( .D(n24765), .E(n6455), .CP(clk), .QN(n5125) );
  EDFD1 \Mem_reg[61][21]  ( .D(n24765), .E(n6454), .CP(clk), .QN(n17990) );
  EDFD1 \Mem_reg[60][21]  ( .D(n24765), .E(n6453), .CP(clk), .QN(n17989) );
  EDFD1 \Mem_reg[59][21]  ( .D(n24765), .E(n6452), .CP(clk), .QN(n4981) );
  EDFD1 \Mem_reg[58][21]  ( .D(n24765), .E(n6451), .CP(clk), .QN(n4933) );
  EDFD1 \Mem_reg[57][21]  ( .D(n24765), .E(n6450), .CP(clk), .QN(n4885) );
  EDFD1 \Mem_reg[56][21]  ( .D(n24765), .E(n6449), .CP(clk), .QN(n4837) );
  EDFD1 \Mem_reg[55][21]  ( .D(n24765), .E(n6448), .CP(clk), .QN(n4789) );
  EDFD1 \Mem_reg[54][21]  ( .D(n24765), .E(n6447), .CP(clk), .QN(n15532) );
  EDFD1 \Mem_reg[53][21]  ( .D(n24765), .E(n6446), .CP(clk), .QN(n4693) );
  EDFD1 \Mem_reg[52][21]  ( .D(n24765), .E(n6445), .CP(clk), .Q(n27120) );
  EDFD1 \Mem_reg[51][21]  ( .D(n24765), .E(n6444), .CP(clk), .QN(n4597) );
  EDFD1 \Mem_reg[50][21]  ( .D(n24765), .E(n6443), .CP(clk), .QN(n4549) );
  EDFD1 \Mem_reg[49][21]  ( .D(n24765), .E(n6442), .CP(clk), .QN(n4501) );
  EDFD1 \Mem_reg[48][21]  ( .D(n24765), .E(n6441), .CP(clk), .QN(n4453) );
  EDFD1 \Mem_reg[47][21]  ( .D(n24765), .E(n6440), .CP(clk), .QN(n4405) );
  EDFD1 \Mem_reg[46][21]  ( .D(n24765), .E(n6439), .CP(clk), .QN(n4357) );
  EDFD1 \Mem_reg[43][21]  ( .D(n24765), .E(n6438), .CP(clk), .QN(n4309) );
  EDFD1 \Mem_reg[42][21]  ( .D(n24765), .E(n6437), .CP(clk), .QN(n4261) );
  EDFD1 \Mem_reg[41][21]  ( .D(n24765), .E(n6436), .CP(clk), .QN(n4213) );
  EDFD1 \Mem_reg[40][21]  ( .D(n24765), .E(n6435), .CP(clk), .QN(n4165) );
  EDFD1 \Mem_reg[39][21]  ( .D(n24765), .E(n6434), .CP(clk), .QN(n4117) );
  EDFD1 \Mem_reg[38][21]  ( .D(n24765), .E(n6433), .CP(clk), .QN(n4069) );
  EDFD1 \Mem_reg[37][21]  ( .D(n24765), .E(n6432), .CP(clk), .QN(n4021) );
  EDFD1 \Mem_reg[36][21]  ( .D(n24765), .E(n6431), .CP(clk), .QN(n3973) );
  EDFD1 \Mem_reg[35][21]  ( .D(n24765), .E(n6430), .CP(clk), .QN(n3925) );
  EDFD1 \Mem_reg[34][21]  ( .D(n24765), .E(n6429), .CP(clk), .QN(n3877) );
  EDFD1 \Mem_reg[33][21]  ( .D(n24765), .E(n6428), .CP(clk), .QN(n3829) );
  EDFD1 \Mem_reg[32][21]  ( .D(n24765), .E(n6427), .CP(clk), .QN(n3781) );
  EDFD1 \Mem_reg[31][21]  ( .D(n24765), .E(n6426), .CP(clk), .QN(n3733) );
  EDFD1 \Mem_reg[30][21]  ( .D(n24765), .E(n6425), .CP(clk), .QN(n3685) );
  EDFD1 \Mem_reg[29][21]  ( .D(n24765), .E(n6424), .CP(clk), .QN(n3637) );
  EDFD1 \Mem_reg[28][21]  ( .D(n24765), .E(n6423), .CP(clk), .QN(n3589) );
  EDFD1 \Mem_reg[27][21]  ( .D(n24765), .E(n6422), .CP(clk), .QN(n3541) );
  EDFD1 \Mem_reg[26][21]  ( .D(n24765), .E(n6421), .CP(clk), .QN(n3493) );
  EDFD1 \Mem_reg[25][21]  ( .D(n24765), .E(n6420), .CP(clk), .QN(n3445) );
  EDFD1 \Mem_reg[24][21]  ( .D(n24765), .E(n6463), .CP(clk), .QN(n3397) );
  EDFD1 \Mem_reg[23][21]  ( .D(n24765), .E(n6464), .CP(clk), .QN(n3349) );
  EDFD1 \Mem_reg[22][21]  ( .D(n24765), .E(n6465), .CP(clk), .QN(n3301) );
  EDFD1 \Mem_reg[21][21]  ( .D(n24765), .E(n6466), .CP(clk), .QN(n3253) );
  EDFD1 \Mem_reg[20][21]  ( .D(n24765), .E(n6467), .CP(clk), .QN(n3205) );
  EDFD1 \Mem_reg[19][21]  ( .D(n24765), .E(n6468), .CP(clk), .QN(n3157) );
  EDFD1 \Mem_reg[18][21]  ( .D(n24765), .E(n6469), .CP(clk), .QN(n3109) );
  EDFD1 \Mem_reg[17][21]  ( .D(n24765), .E(n6470), .CP(clk), .QN(n3061) );
  EDFD1 \Mem_reg[16][21]  ( .D(n24765), .E(n6471), .CP(clk), .QN(n3013) );
  EDFD1 \Mem_reg[15][21]  ( .D(n24765), .E(n6472), .CP(clk), .QN(n2965) );
  EDFD1 \Mem_reg[14][21]  ( .D(n24765), .E(n24720), .CP(clk), .QN(n2917) );
  EDFD1 \Mem_reg[13][21]  ( .D(n24765), .E(n24709), .CP(clk), .QN(n2869) );
  EDFD1 \Mem_reg[12][21]  ( .D(n24765), .E(n24717), .CP(clk), .QN(n2821) );
  EDFD1 \Mem_reg[11][21]  ( .D(n24765), .E(n24707), .CP(clk), .QN(n2773) );
  EDFD1 \Mem_reg[10][21]  ( .D(n24765), .E(n6477), .CP(clk), .QN(n2725) );
  EDFD1 \Mem_reg[9][21]  ( .D(n24765), .E(n24708), .CP(clk), .QN(n2677) );
  EDFD1 \Mem_reg[8][21]  ( .D(n24765), .E(n15642), .CP(clk), .QN(n2629) );
  EDFD1 \Mem_reg[7][21]  ( .D(n24765), .E(n24718), .CP(clk), .QN(n2581) );
  EDFD1 \Mem_reg[6][21]  ( .D(n24765), .E(n24716), .CP(clk), .QN(n2533) );
  EDFD1 \Mem_reg[5][21]  ( .D(n24765), .E(n24719), .CP(clk), .QN(n2485) );
  EDFD1 \Mem_reg[4][21]  ( .D(n24765), .E(n24706), .CP(clk), .QN(n2437) );
  EDFD1 \Mem_reg[3][21]  ( .D(n24765), .E(n24721), .CP(clk), .QN(n2389) );
  EDFD1 \Mem_reg[2][21]  ( .D(n24765), .E(n6460), .CP(clk), .QN(n2341) );
  EDFD1 \Mem_reg[1][21]  ( .D(n24765), .E(n24703), .CP(clk), .QN(n2293) );
  EDFD1 \Mem_reg[0][21]  ( .D(n24765), .E(n24705), .CP(clk), .QN(n2245) );
  EDFD1 \Mem_reg[88][20]  ( .D(n24763), .E(n6419), .CP(clk), .Q(n27117) );
  EDFD1 \Mem_reg[87][20]  ( .D(n24763), .E(n6418), .CP(clk), .QN(n6326) );
  EDFD1 \Mem_reg[86][20]  ( .D(n24763), .E(n6417), .CP(clk), .QN(n24619) );
  EDFD1 \Mem_reg[85][20]  ( .D(n24763), .E(n6416), .CP(clk), .QN(n6230) );
  EDFD1 \Mem_reg[84][20]  ( .D(n24763), .E(n6415), .CP(clk), .QN(n6182) );
  EDFD1 \Mem_reg[83][20]  ( .D(n24763), .E(n6414), .CP(clk), .QN(n6134) );
  EDFD1 \Mem_reg[82][20]  ( .D(n24763), .E(n6413), .CP(clk), .QN(n6086) );
  EDFD1 \Mem_reg[81][20]  ( .D(n24763), .E(n6412), .CP(clk), .QN(n6038) );
  EDFD1 \Mem_reg[80][20]  ( .D(n24763), .E(n6411), .CP(clk), .QN(n5990) );
  EDFD1 \Mem_reg[79][20]  ( .D(n24763), .E(n6410), .CP(clk), .QN(n5942) );
  EDFD1 \Mem_reg[78][20]  ( .D(n24763), .E(n6409), .CP(clk), .QN(n5894) );
  EDFD1 \Mem_reg[77][20]  ( .D(n24763), .E(n6408), .CP(clk), .QN(n5846) );
  EDFD1 \Mem_reg[76][20]  ( .D(n24763), .E(n6407), .CP(clk), .QN(n5798) );
  EDFD1 \Mem_reg[75][20]  ( .D(n24763), .E(n6406), .CP(clk), .QN(n27118) );
  EDFD1 \Mem_reg[74][20]  ( .D(n24763), .E(n6405), .CP(clk), .QN(n5702) );
  EDFD1 \Mem_reg[73][20]  ( .D(n24763), .E(n6404), .CP(clk), .QN(n27119) );
  EDFD1 \Mem_reg[72][20]  ( .D(n24763), .E(n6403), .CP(clk), .QN(n5606) );
  EDFD1 \Mem_reg[71][20]  ( .D(n24763), .E(n6402), .CP(clk), .QN(n5558) );
  EDFD1 \Mem_reg[70][20]  ( .D(n24763), .E(n6401), .CP(clk), .QN(n5510) );
  EDFD1 \Mem_reg[69][20]  ( .D(n24763), .E(n6400), .CP(clk), .QN(n5462) );
  EDFD1 \Mem_reg[68][20]  ( .D(n24763), .E(n6399), .CP(clk), .QN(n5414) );
  EDFD1 \Mem_reg[67][20]  ( .D(n24763), .E(n6398), .CP(clk), .QN(n5366) );
  EDFD1 \Mem_reg[66][20]  ( .D(n24763), .E(n6397), .CP(clk), .QN(n5318) );
  EDFD1 \Mem_reg[65][20]  ( .D(n24763), .E(n6396), .CP(clk), .QN(n15529) );
  EDFD1 \Mem_reg[64][20]  ( .D(n24763), .E(n6395), .CP(clk), .QN(n5222) );
  EDFD1 \Mem_reg[63][20]  ( .D(n24763), .E(n6456), .CP(clk), .QN(n5174) );
  EDFD1 \Mem_reg[62][20]  ( .D(n24763), .E(n6455), .CP(clk), .QN(n5126) );
  EDFD1 \Mem_reg[61][20]  ( .D(n24763), .E(n6454), .CP(clk), .QN(n17987) );
  EDFD1 \Mem_reg[60][20]  ( .D(n24763), .E(n6453), .CP(clk), .QN(n17986) );
  EDFD1 \Mem_reg[59][20]  ( .D(n24763), .E(n6452), .CP(clk), .QN(n4982) );
  EDFD1 \Mem_reg[58][20]  ( .D(n24763), .E(n6451), .CP(clk), .QN(n4934) );
  EDFD1 \Mem_reg[57][20]  ( .D(n24763), .E(n6450), .CP(clk), .QN(n4886) );
  EDFD1 \Mem_reg[56][20]  ( .D(n24763), .E(n6449), .CP(clk), .QN(n4838) );
  EDFD1 \Mem_reg[55][20]  ( .D(n24763), .E(n6448), .CP(clk), .QN(n4790) );
  EDFD1 \Mem_reg[54][20]  ( .D(n24763), .E(n6447), .CP(clk), .QN(n15528) );
  EDFD1 \Mem_reg[53][20]  ( .D(n24763), .E(n6446), .CP(clk), .QN(n4694) );
  EDFD1 \Mem_reg[52][20]  ( .D(n24763), .E(n6445), .CP(clk), .Q(n27116) );
  EDFD1 \Mem_reg[51][20]  ( .D(n24763), .E(n6444), .CP(clk), .QN(n4598) );
  EDFD1 \Mem_reg[50][20]  ( .D(n24763), .E(n6443), .CP(clk), .QN(n4550) );
  EDFD1 \Mem_reg[49][20]  ( .D(n24763), .E(n6442), .CP(clk), .QN(n4502) );
  EDFD1 \Mem_reg[48][20]  ( .D(n24763), .E(n6441), .CP(clk), .QN(n4454) );
  EDFD1 \Mem_reg[47][20]  ( .D(n24763), .E(n6440), .CP(clk), .QN(n4406) );
  EDFD1 \Mem_reg[46][20]  ( .D(n24763), .E(n6439), .CP(clk), .QN(n4358) );
  EDFD1 \Mem_reg[43][20]  ( .D(n24763), .E(n6438), .CP(clk), .QN(n4310) );
  EDFD1 \Mem_reg[42][20]  ( .D(n24763), .E(n6437), .CP(clk), .QN(n4262) );
  EDFD1 \Mem_reg[41][20]  ( .D(n24763), .E(n6436), .CP(clk), .QN(n4214) );
  EDFD1 \Mem_reg[40][20]  ( .D(n24763), .E(n6435), .CP(clk), .QN(n4166) );
  EDFD1 \Mem_reg[39][20]  ( .D(n24763), .E(n6434), .CP(clk), .QN(n4118) );
  EDFD1 \Mem_reg[38][20]  ( .D(n24763), .E(n6433), .CP(clk), .QN(n4070) );
  EDFD1 \Mem_reg[37][20]  ( .D(n24763), .E(n6432), .CP(clk), .QN(n4022) );
  EDFD1 \Mem_reg[36][20]  ( .D(n24763), .E(n6431), .CP(clk), .QN(n3974) );
  EDFD1 \Mem_reg[35][20]  ( .D(n24763), .E(n6430), .CP(clk), .QN(n3926) );
  EDFD1 \Mem_reg[34][20]  ( .D(n24763), .E(n6429), .CP(clk), .QN(n3878) );
  EDFD1 \Mem_reg[33][20]  ( .D(n24763), .E(n6428), .CP(clk), .QN(n3830) );
  EDFD1 \Mem_reg[32][20]  ( .D(n24763), .E(n6427), .CP(clk), .QN(n3782) );
  EDFD1 \Mem_reg[31][20]  ( .D(n24763), .E(n6426), .CP(clk), .QN(n3734) );
  EDFD1 \Mem_reg[30][20]  ( .D(n24763), .E(n6425), .CP(clk), .QN(n3686) );
  EDFD1 \Mem_reg[29][20]  ( .D(n24763), .E(n6424), .CP(clk), .QN(n3638) );
  EDFD1 \Mem_reg[28][20]  ( .D(n24763), .E(n6423), .CP(clk), .QN(n3590) );
  EDFD1 \Mem_reg[27][20]  ( .D(n24763), .E(n6422), .CP(clk), .QN(n3542) );
  EDFD1 \Mem_reg[26][20]  ( .D(n24763), .E(n6421), .CP(clk), .QN(n3494) );
  EDFD1 \Mem_reg[25][20]  ( .D(n24763), .E(n6420), .CP(clk), .QN(n3446) );
  EDFD1 \Mem_reg[24][20]  ( .D(n24763), .E(n6463), .CP(clk), .QN(n3398) );
  EDFD1 \Mem_reg[23][20]  ( .D(n24763), .E(n6464), .CP(clk), .QN(n3350) );
  EDFD1 \Mem_reg[22][20]  ( .D(n24763), .E(n6465), .CP(clk), .QN(n3302) );
  EDFD1 \Mem_reg[21][20]  ( .D(n24763), .E(n6466), .CP(clk), .QN(n3254) );
  EDFD1 \Mem_reg[20][20]  ( .D(n24763), .E(n6467), .CP(clk), .QN(n3206) );
  EDFD1 \Mem_reg[19][20]  ( .D(n24763), .E(n6468), .CP(clk), .QN(n3158) );
  EDFD1 \Mem_reg[18][20]  ( .D(n24763), .E(n6469), .CP(clk), .QN(n3110) );
  EDFD1 \Mem_reg[17][20]  ( .D(n24763), .E(n6470), .CP(clk), .QN(n3062) );
  EDFD1 \Mem_reg[16][20]  ( .D(n24763), .E(n6471), .CP(clk), .QN(n3014) );
  EDFD1 \Mem_reg[15][20]  ( .D(n24763), .E(n6472), .CP(clk), .QN(n2966) );
  EDFD1 \Mem_reg[14][20]  ( .D(n24763), .E(n24720), .CP(clk), .QN(n2918) );
  EDFD1 \Mem_reg[13][20]  ( .D(n24763), .E(n24709), .CP(clk), .QN(n2870) );
  EDFD1 \Mem_reg[12][20]  ( .D(n24763), .E(n24717), .CP(clk), .QN(n2822) );
  EDFD1 \Mem_reg[11][20]  ( .D(n24763), .E(n24707), .CP(clk), .QN(n2774) );
  EDFD1 \Mem_reg[10][20]  ( .D(n24763), .E(n6477), .CP(clk), .QN(n2726) );
  EDFD1 \Mem_reg[9][20]  ( .D(n24763), .E(n24708), .CP(clk), .QN(n2678) );
  EDFD1 \Mem_reg[8][20]  ( .D(n24763), .E(n15642), .CP(clk), .QN(n2630) );
  EDFD1 \Mem_reg[7][20]  ( .D(n24763), .E(n24718), .CP(clk), .QN(n2582) );
  EDFD1 \Mem_reg[6][20]  ( .D(n24763), .E(n24716), .CP(clk), .QN(n2534) );
  EDFD1 \Mem_reg[5][20]  ( .D(n24763), .E(n24719), .CP(clk), .QN(n2486) );
  EDFD1 \Mem_reg[4][20]  ( .D(n24763), .E(n24706), .CP(clk), .QN(n2438) );
  EDFD1 \Mem_reg[3][20]  ( .D(n24763), .E(n24721), .CP(clk), .QN(n2390) );
  EDFD1 \Mem_reg[2][20]  ( .D(n24763), .E(n6460), .CP(clk), .QN(n2342) );
  EDFD1 \Mem_reg[1][20]  ( .D(n24763), .E(n24703), .CP(clk), .QN(n2294) );
  EDFD1 \Mem_reg[0][20]  ( .D(n24763), .E(n24705), .CP(clk), .QN(n2246) );
  EDFD1 \Mem_reg[88][19]  ( .D(n24761), .E(n6419), .CP(clk), .Q(n27113) );
  EDFD1 \Mem_reg[5][19]  ( .D(n24761), .E(n24719), .CP(clk), .QN(n2487) );
  EDFD1 \Mem_reg[4][19]  ( .D(n24761), .E(n24706), .CP(clk), .QN(n2439) );
  EDFD1 \Mem_reg[3][19]  ( .D(n24761), .E(n24721), .CP(clk), .QN(n2391) );
  EDFD1 \Mem_reg[2][19]  ( .D(n24761), .E(n6460), .CP(clk), .QN(n2343) );
  EDFD1 \Mem_reg[1][19]  ( .D(n24761), .E(n24703), .CP(clk), .QN(n2295) );
  EDFD1 \Mem_reg[0][19]  ( .D(n24761), .E(n24705), .CP(clk), .QN(n2247) );
  EDFD1 \Mem_reg[87][19]  ( .D(n24761), .E(n6418), .CP(clk), .QN(n6327) );
  EDFD1 \Mem_reg[86][19]  ( .D(n24761), .E(n6417), .CP(clk), .QN(n24616) );
  EDFD1 \Mem_reg[85][19]  ( .D(n24761), .E(n6416), .CP(clk), .QN(n6231) );
  EDFD1 \Mem_reg[84][19]  ( .D(n24761), .E(n6415), .CP(clk), .QN(n6183) );
  EDFD1 \Mem_reg[83][19]  ( .D(n24761), .E(n6414), .CP(clk), .QN(n6135) );
  EDFD1 \Mem_reg[82][19]  ( .D(n24761), .E(n6413), .CP(clk), .QN(n6087) );
  EDFD1 \Mem_reg[81][19]  ( .D(n24761), .E(n6412), .CP(clk), .QN(n6039) );
  EDFD1 \Mem_reg[80][19]  ( .D(n24761), .E(n6411), .CP(clk), .QN(n5991) );
  EDFD1 \Mem_reg[79][19]  ( .D(n24761), .E(n6410), .CP(clk), .QN(n5943) );
  EDFD1 \Mem_reg[78][19]  ( .D(n24761), .E(n6409), .CP(clk), .QN(n5895) );
  EDFD1 \Mem_reg[77][19]  ( .D(n24761), .E(n6408), .CP(clk), .QN(n5847) );
  EDFD1 \Mem_reg[76][19]  ( .D(n24761), .E(n6407), .CP(clk), .QN(n5799) );
  EDFD1 \Mem_reg[75][19]  ( .D(n24761), .E(n6406), .CP(clk), .QN(n27114) );
  EDFD1 \Mem_reg[74][19]  ( .D(n24761), .E(n6405), .CP(clk), .QN(n5703) );
  EDFD1 \Mem_reg[73][19]  ( .D(n24761), .E(n6404), .CP(clk), .QN(n27115) );
  EDFD1 \Mem_reg[72][19]  ( .D(n24761), .E(n6403), .CP(clk), .QN(n5607) );
  EDFD1 \Mem_reg[71][19]  ( .D(n24761), .E(n6402), .CP(clk), .QN(n5559) );
  EDFD1 \Mem_reg[70][19]  ( .D(n24761), .E(n6401), .CP(clk), .QN(n5511) );
  EDFD1 \Mem_reg[69][19]  ( .D(n24761), .E(n6400), .CP(clk), .QN(n5463) );
  EDFD1 \Mem_reg[68][19]  ( .D(n24761), .E(n6399), .CP(clk), .QN(n5415) );
  EDFD1 \Mem_reg[67][19]  ( .D(n24761), .E(n6398), .CP(clk), .QN(n5367) );
  EDFD1 \Mem_reg[66][19]  ( .D(n24761), .E(n6397), .CP(clk), .QN(n5319) );
  EDFD1 \Mem_reg[65][19]  ( .D(n24761), .E(n6396), .CP(clk), .QN(n15525) );
  EDFD1 \Mem_reg[64][19]  ( .D(n24761), .E(n6395), .CP(clk), .QN(n5223) );
  EDFD1 \Mem_reg[63][19]  ( .D(n24761), .E(n6456), .CP(clk), .QN(n5175) );
  EDFD1 \Mem_reg[62][19]  ( .D(n24761), .E(n6455), .CP(clk), .QN(n5127) );
  EDFD1 \Mem_reg[61][19]  ( .D(n24761), .E(n6454), .CP(clk), .QN(n17984) );
  EDFD1 \Mem_reg[60][19]  ( .D(n24761), .E(n6453), .CP(clk), .QN(n17983) );
  EDFD1 \Mem_reg[59][19]  ( .D(n24761), .E(n6452), .CP(clk), .QN(n4983) );
  EDFD1 \Mem_reg[58][19]  ( .D(n24761), .E(n6451), .CP(clk), .QN(n4935) );
  EDFD1 \Mem_reg[57][19]  ( .D(n24761), .E(n6450), .CP(clk), .QN(n4887) );
  EDFD1 \Mem_reg[56][19]  ( .D(n24761), .E(n6449), .CP(clk), .QN(n4839) );
  EDFD1 \Mem_reg[55][19]  ( .D(n24761), .E(n6448), .CP(clk), .QN(n4791) );
  EDFD1 \Mem_reg[54][19]  ( .D(n24761), .E(n6447), .CP(clk), .QN(n15524) );
  EDFD1 \Mem_reg[53][19]  ( .D(n24761), .E(n6446), .CP(clk), .QN(n4695) );
  EDFD1 \Mem_reg[52][19]  ( .D(n24761), .E(n6445), .CP(clk), .Q(n27112) );
  EDFD1 \Mem_reg[51][19]  ( .D(n24761), .E(n6444), .CP(clk), .QN(n4599) );
  EDFD1 \Mem_reg[50][19]  ( .D(n24761), .E(n6443), .CP(clk), .QN(n4551) );
  EDFD1 \Mem_reg[49][19]  ( .D(n24761), .E(n6442), .CP(clk), .QN(n4503) );
  EDFD1 \Mem_reg[48][19]  ( .D(n24761), .E(n6441), .CP(clk), .QN(n4455) );
  EDFD1 \Mem_reg[47][19]  ( .D(n24761), .E(n6440), .CP(clk), .QN(n4407) );
  EDFD1 \Mem_reg[46][19]  ( .D(n24761), .E(n6439), .CP(clk), .QN(n4359) );
  EDFD1 \Mem_reg[43][19]  ( .D(n24761), .E(n6438), .CP(clk), .QN(n4311) );
  EDFD1 \Mem_reg[42][19]  ( .D(n24761), .E(n6437), .CP(clk), .QN(n4263) );
  EDFD1 \Mem_reg[41][19]  ( .D(n24761), .E(n6436), .CP(clk), .QN(n4215) );
  EDFD1 \Mem_reg[40][19]  ( .D(n24761), .E(n6435), .CP(clk), .QN(n4167) );
  EDFD1 \Mem_reg[39][19]  ( .D(n24761), .E(n6434), .CP(clk), .QN(n4119) );
  EDFD1 \Mem_reg[38][19]  ( .D(n24761), .E(n6433), .CP(clk), .QN(n4071) );
  EDFD1 \Mem_reg[37][19]  ( .D(n24761), .E(n6432), .CP(clk), .QN(n4023) );
  EDFD1 \Mem_reg[36][19]  ( .D(n24761), .E(n6431), .CP(clk), .QN(n3975) );
  EDFD1 \Mem_reg[35][19]  ( .D(n24761), .E(n6430), .CP(clk), .QN(n3927) );
  EDFD1 \Mem_reg[34][19]  ( .D(n24761), .E(n6429), .CP(clk), .QN(n3879) );
  EDFD1 \Mem_reg[33][19]  ( .D(n24761), .E(n6428), .CP(clk), .QN(n3831) );
  EDFD1 \Mem_reg[32][19]  ( .D(n24761), .E(n6427), .CP(clk), .QN(n3783) );
  EDFD1 \Mem_reg[31][19]  ( .D(n24761), .E(n6426), .CP(clk), .QN(n3735) );
  EDFD1 \Mem_reg[30][19]  ( .D(n24761), .E(n6425), .CP(clk), .QN(n3687) );
  EDFD1 \Mem_reg[29][19]  ( .D(n24761), .E(n6424), .CP(clk), .QN(n3639) );
  EDFD1 \Mem_reg[28][19]  ( .D(n24761), .E(n6423), .CP(clk), .QN(n3591) );
  EDFD1 \Mem_reg[27][19]  ( .D(n24761), .E(n6422), .CP(clk), .QN(n3543) );
  EDFD1 \Mem_reg[26][19]  ( .D(n24761), .E(n6421), .CP(clk), .QN(n3495) );
  EDFD1 \Mem_reg[25][19]  ( .D(n24761), .E(n6420), .CP(clk), .QN(n3447) );
  EDFD1 \Mem_reg[24][19]  ( .D(n24761), .E(n6463), .CP(clk), .QN(n3399) );
  EDFD1 \Mem_reg[23][19]  ( .D(n24761), .E(n6464), .CP(clk), .QN(n3351) );
  EDFD1 \Mem_reg[22][19]  ( .D(n24761), .E(n6465), .CP(clk), .QN(n3303) );
  EDFD1 \Mem_reg[21][19]  ( .D(n24761), .E(n6466), .CP(clk), .QN(n3255) );
  EDFD1 \Mem_reg[20][19]  ( .D(n24761), .E(n6467), .CP(clk), .QN(n3207) );
  EDFD1 \Mem_reg[19][19]  ( .D(n24761), .E(n6468), .CP(clk), .QN(n3159) );
  EDFD1 \Mem_reg[18][19]  ( .D(n24761), .E(n6469), .CP(clk), .QN(n3111) );
  EDFD1 \Mem_reg[17][19]  ( .D(n24761), .E(n6470), .CP(clk), .QN(n3063) );
  EDFD1 \Mem_reg[16][19]  ( .D(n24761), .E(n6471), .CP(clk), .QN(n3015) );
  EDFD1 \Mem_reg[15][19]  ( .D(n24761), .E(n6472), .CP(clk), .QN(n2967) );
  EDFD1 \Mem_reg[14][19]  ( .D(n24761), .E(n24720), .CP(clk), .QN(n2919) );
  EDFD1 \Mem_reg[13][19]  ( .D(n24761), .E(n24709), .CP(clk), .QN(n2871) );
  EDFD1 \Mem_reg[12][19]  ( .D(n24761), .E(n24717), .CP(clk), .QN(n2823) );
  EDFD1 \Mem_reg[11][19]  ( .D(n24761), .E(n24707), .CP(clk), .QN(n2775) );
  EDFD1 \Mem_reg[10][19]  ( .D(n24761), .E(n6477), .CP(clk), .QN(n2727) );
  EDFD1 \Mem_reg[9][19]  ( .D(n24761), .E(n24708), .CP(clk), .QN(n2679) );
  EDFD1 \Mem_reg[8][19]  ( .D(n24761), .E(n15642), .CP(clk), .QN(n2631) );
  EDFD1 \Mem_reg[7][19]  ( .D(n24761), .E(n24718), .CP(clk), .QN(n2583) );
  EDFD1 \Mem_reg[6][19]  ( .D(n24761), .E(n24716), .CP(clk), .QN(n2535) );
  EDFD1 \Mem_reg[88][18]  ( .D(n24759), .E(n6419), .CP(clk), .Q(n27109) );
  EDFD1 \Mem_reg[87][18]  ( .D(n24759), .E(n6418), .CP(clk), .QN(n6328) );
  EDFD1 \Mem_reg[86][18]  ( .D(n24759), .E(n6417), .CP(clk), .QN(n24613) );
  EDFD1 \Mem_reg[85][18]  ( .D(n24759), .E(n6416), .CP(clk), .QN(n6232) );
  EDFD1 \Mem_reg[84][18]  ( .D(n24759), .E(n6415), .CP(clk), .QN(n6184) );
  EDFD1 \Mem_reg[83][18]  ( .D(n24759), .E(n6414), .CP(clk), .QN(n6136) );
  EDFD1 \Mem_reg[82][18]  ( .D(n24759), .E(n6413), .CP(clk), .QN(n6088) );
  EDFD1 \Mem_reg[81][18]  ( .D(n24759), .E(n6412), .CP(clk), .QN(n6040) );
  EDFD1 \Mem_reg[80][18]  ( .D(n24759), .E(n6411), .CP(clk), .QN(n5992) );
  EDFD1 \Mem_reg[79][18]  ( .D(n24759), .E(n6410), .CP(clk), .QN(n5944) );
  EDFD1 \Mem_reg[78][18]  ( .D(n24759), .E(n6409), .CP(clk), .QN(n5896) );
  EDFD1 \Mem_reg[77][18]  ( .D(n24759), .E(n6408), .CP(clk), .QN(n5848) );
  EDFD1 \Mem_reg[76][18]  ( .D(n24759), .E(n6407), .CP(clk), .QN(n5800) );
  EDFD1 \Mem_reg[75][18]  ( .D(n24759), .E(n6406), .CP(clk), .QN(n27110) );
  EDFD1 \Mem_reg[74][18]  ( .D(n24759), .E(n6405), .CP(clk), .QN(n5704) );
  EDFD1 \Mem_reg[73][18]  ( .D(n24759), .E(n6404), .CP(clk), .QN(n27111) );
  EDFD1 \Mem_reg[72][18]  ( .D(n24759), .E(n6403), .CP(clk), .QN(n5608) );
  EDFD1 \Mem_reg[71][18]  ( .D(n24759), .E(n6402), .CP(clk), .QN(n5560) );
  EDFD1 \Mem_reg[70][18]  ( .D(n24759), .E(n6401), .CP(clk), .QN(n5512) );
  EDFD1 \Mem_reg[69][18]  ( .D(n24759), .E(n6400), .CP(clk), .QN(n5464) );
  EDFD1 \Mem_reg[68][18]  ( .D(n24759), .E(n6399), .CP(clk), .QN(n5416) );
  EDFD1 \Mem_reg[67][18]  ( .D(n24759), .E(n6398), .CP(clk), .QN(n5368) );
  EDFD1 \Mem_reg[66][18]  ( .D(n24759), .E(n6397), .CP(clk), .QN(n5320) );
  EDFD1 \Mem_reg[65][18]  ( .D(n24759), .E(n6396), .CP(clk), .QN(n15521) );
  EDFD1 \Mem_reg[64][18]  ( .D(n24759), .E(n6395), .CP(clk), .QN(n5224) );
  EDFD1 \Mem_reg[63][18]  ( .D(n24759), .E(n6456), .CP(clk), .QN(n5176) );
  EDFD1 \Mem_reg[62][18]  ( .D(n24759), .E(n6455), .CP(clk), .QN(n5128) );
  EDFD1 \Mem_reg[61][18]  ( .D(n24759), .E(n6454), .CP(clk), .QN(n17981) );
  EDFD1 \Mem_reg[60][18]  ( .D(n24759), .E(n6453), .CP(clk), .QN(n17980) );
  EDFD1 \Mem_reg[59][18]  ( .D(n24759), .E(n6452), .CP(clk), .QN(n4984) );
  EDFD1 \Mem_reg[58][18]  ( .D(n24759), .E(n6451), .CP(clk), .QN(n4936) );
  EDFD1 \Mem_reg[57][18]  ( .D(n24759), .E(n6450), .CP(clk), .QN(n4888) );
  EDFD1 \Mem_reg[56][18]  ( .D(n24759), .E(n6449), .CP(clk), .QN(n4840) );
  EDFD1 \Mem_reg[55][18]  ( .D(n24759), .E(n6448), .CP(clk), .QN(n4792) );
  EDFD1 \Mem_reg[54][18]  ( .D(n24759), .E(n6447), .CP(clk), .QN(n15520) );
  EDFD1 \Mem_reg[53][18]  ( .D(n24759), .E(n6446), .CP(clk), .QN(n4696) );
  EDFD1 \Mem_reg[52][18]  ( .D(n24759), .E(n6445), .CP(clk), .Q(n27108) );
  EDFD1 \Mem_reg[51][18]  ( .D(n24759), .E(n6444), .CP(clk), .QN(n4600) );
  EDFD1 \Mem_reg[50][18]  ( .D(n24759), .E(n6443), .CP(clk), .QN(n4552) );
  EDFD1 \Mem_reg[49][18]  ( .D(n24759), .E(n6442), .CP(clk), .QN(n4504) );
  EDFD1 \Mem_reg[48][18]  ( .D(n24759), .E(n6441), .CP(clk), .QN(n4456) );
  EDFD1 \Mem_reg[47][18]  ( .D(n24759), .E(n6440), .CP(clk), .QN(n4408) );
  EDFD1 \Mem_reg[46][18]  ( .D(n24759), .E(n6439), .CP(clk), .QN(n4360) );
  EDFD1 \Mem_reg[43][18]  ( .D(n24759), .E(n6438), .CP(clk), .QN(n4312) );
  EDFD1 \Mem_reg[42][18]  ( .D(n24759), .E(n6437), .CP(clk), .QN(n4264) );
  EDFD1 \Mem_reg[41][18]  ( .D(n24759), .E(n6436), .CP(clk), .QN(n4216) );
  EDFD1 \Mem_reg[40][18]  ( .D(n24759), .E(n6435), .CP(clk), .QN(n4168) );
  EDFD1 \Mem_reg[39][18]  ( .D(n24759), .E(n6434), .CP(clk), .QN(n4120) );
  EDFD1 \Mem_reg[38][18]  ( .D(n24759), .E(n6433), .CP(clk), .QN(n4072) );
  EDFD1 \Mem_reg[37][18]  ( .D(n24759), .E(n6432), .CP(clk), .QN(n4024) );
  EDFD1 \Mem_reg[36][18]  ( .D(n24759), .E(n6431), .CP(clk), .QN(n3976) );
  EDFD1 \Mem_reg[35][18]  ( .D(n24759), .E(n6430), .CP(clk), .QN(n3928) );
  EDFD1 \Mem_reg[34][18]  ( .D(n24759), .E(n6429), .CP(clk), .QN(n3880) );
  EDFD1 \Mem_reg[33][18]  ( .D(n24759), .E(n6428), .CP(clk), .QN(n3832) );
  EDFD1 \Mem_reg[32][18]  ( .D(n24759), .E(n6427), .CP(clk), .QN(n3784) );
  EDFD1 \Mem_reg[31][18]  ( .D(n24759), .E(n6426), .CP(clk), .QN(n3736) );
  EDFD1 \Mem_reg[30][18]  ( .D(n24759), .E(n6425), .CP(clk), .QN(n3688) );
  EDFD1 \Mem_reg[29][18]  ( .D(n24759), .E(n6424), .CP(clk), .QN(n3640) );
  EDFD1 \Mem_reg[28][18]  ( .D(n24759), .E(n6423), .CP(clk), .QN(n3592) );
  EDFD1 \Mem_reg[27][18]  ( .D(n24759), .E(n6422), .CP(clk), .QN(n3544) );
  EDFD1 \Mem_reg[26][18]  ( .D(n24759), .E(n6421), .CP(clk), .QN(n3496) );
  EDFD1 \Mem_reg[25][18]  ( .D(n24759), .E(n6420), .CP(clk), .QN(n3448) );
  EDFD1 \Mem_reg[24][18]  ( .D(n24759), .E(n6463), .CP(clk), .QN(n3400) );
  EDFD1 \Mem_reg[23][18]  ( .D(n24759), .E(n6464), .CP(clk), .QN(n3352) );
  EDFD1 \Mem_reg[22][18]  ( .D(n24759), .E(n6465), .CP(clk), .QN(n3304) );
  EDFD1 \Mem_reg[21][18]  ( .D(n24759), .E(n6466), .CP(clk), .QN(n3256) );
  EDFD1 \Mem_reg[20][18]  ( .D(n24759), .E(n6467), .CP(clk), .QN(n3208) );
  EDFD1 \Mem_reg[19][18]  ( .D(n24759), .E(n6468), .CP(clk), .QN(n3160) );
  EDFD1 \Mem_reg[18][18]  ( .D(n24759), .E(n6469), .CP(clk), .QN(n3112) );
  EDFD1 \Mem_reg[17][18]  ( .D(n24759), .E(n6470), .CP(clk), .QN(n3064) );
  EDFD1 \Mem_reg[16][18]  ( .D(n24759), .E(n6471), .CP(clk), .QN(n3016) );
  EDFD1 \Mem_reg[15][18]  ( .D(n24759), .E(n6472), .CP(clk), .QN(n2968) );
  EDFD1 \Mem_reg[14][18]  ( .D(n24759), .E(n24720), .CP(clk), .QN(n2920) );
  EDFD1 \Mem_reg[13][18]  ( .D(n24759), .E(n24709), .CP(clk), .QN(n2872) );
  EDFD1 \Mem_reg[12][18]  ( .D(n24759), .E(n24717), .CP(clk), .QN(n2824) );
  EDFD1 \Mem_reg[11][18]  ( .D(n24759), .E(n24707), .CP(clk), .QN(n2776) );
  EDFD1 \Mem_reg[10][18]  ( .D(n24759), .E(n6477), .CP(clk), .QN(n2728) );
  EDFD1 \Mem_reg[9][18]  ( .D(n24759), .E(n24708), .CP(clk), .QN(n2680) );
  EDFD1 \Mem_reg[8][18]  ( .D(n24759), .E(n15642), .CP(clk), .QN(n2632) );
  EDFD1 \Mem_reg[7][18]  ( .D(n24759), .E(n24718), .CP(clk), .QN(n2584) );
  EDFD1 \Mem_reg[6][18]  ( .D(n24759), .E(n24716), .CP(clk), .QN(n2536) );
  EDFD1 \Mem_reg[5][18]  ( .D(n24759), .E(n24719), .CP(clk), .QN(n2488) );
  EDFD1 \Mem_reg[4][18]  ( .D(n24759), .E(n24706), .CP(clk), .QN(n2440) );
  EDFD1 \Mem_reg[3][18]  ( .D(n24759), .E(n24721), .CP(clk), .QN(n2392) );
  EDFD1 \Mem_reg[2][18]  ( .D(n24759), .E(n6460), .CP(clk), .QN(n2344) );
  EDFD1 \Mem_reg[1][18]  ( .D(n24759), .E(n24703), .CP(clk), .QN(n2296) );
  EDFD1 \Mem_reg[0][18]  ( .D(n24759), .E(n24705), .CP(clk), .QN(n2248) );
  EDFD1 \Mem_reg[88][17]  ( .D(n24757), .E(n6419), .CP(clk), .Q(n27105) );
  EDFD1 \Mem_reg[87][17]  ( .D(n24757), .E(n6418), .CP(clk), .QN(n6329) );
  EDFD1 \Mem_reg[86][17]  ( .D(n24757), .E(n6417), .CP(clk), .QN(n24610) );
  EDFD1 \Mem_reg[85][17]  ( .D(n24757), .E(n6416), .CP(clk), .QN(n6233) );
  EDFD1 \Mem_reg[84][17]  ( .D(n24757), .E(n6415), .CP(clk), .QN(n6185) );
  EDFD1 \Mem_reg[83][17]  ( .D(n24757), .E(n6414), .CP(clk), .QN(n6137) );
  EDFD1 \Mem_reg[82][17]  ( .D(n24757), .E(n6413), .CP(clk), .QN(n6089) );
  EDFD1 \Mem_reg[81][17]  ( .D(n24757), .E(n6412), .CP(clk), .QN(n6041) );
  EDFD1 \Mem_reg[80][17]  ( .D(n24757), .E(n6411), .CP(clk), .QN(n5993) );
  EDFD1 \Mem_reg[79][17]  ( .D(n24757), .E(n6410), .CP(clk), .QN(n5945) );
  EDFD1 \Mem_reg[78][17]  ( .D(n24757), .E(n6409), .CP(clk), .QN(n5897) );
  EDFD1 \Mem_reg[77][17]  ( .D(n24757), .E(n6408), .CP(clk), .QN(n5849) );
  EDFD1 \Mem_reg[76][17]  ( .D(n24757), .E(n6407), .CP(clk), .QN(n5801) );
  EDFD1 \Mem_reg[75][17]  ( .D(n24757), .E(n6406), .CP(clk), .QN(n27106) );
  EDFD1 \Mem_reg[74][17]  ( .D(n24757), .E(n6405), .CP(clk), .QN(n5705) );
  EDFD1 \Mem_reg[73][17]  ( .D(n24757), .E(n6404), .CP(clk), .QN(n27107) );
  EDFD1 \Mem_reg[72][17]  ( .D(n24757), .E(n6403), .CP(clk), .QN(n5609) );
  EDFD1 \Mem_reg[71][17]  ( .D(n24757), .E(n6402), .CP(clk), .QN(n5561) );
  EDFD1 \Mem_reg[70][17]  ( .D(n24757), .E(n6401), .CP(clk), .QN(n5513) );
  EDFD1 \Mem_reg[69][17]  ( .D(n24757), .E(n6400), .CP(clk), .QN(n5465) );
  EDFD1 \Mem_reg[68][17]  ( .D(n24757), .E(n6399), .CP(clk), .QN(n5417) );
  EDFD1 \Mem_reg[67][17]  ( .D(n24757), .E(n6398), .CP(clk), .QN(n5369) );
  EDFD1 \Mem_reg[66][17]  ( .D(n24757), .E(n6397), .CP(clk), .QN(n5321) );
  EDFD1 \Mem_reg[65][17]  ( .D(n24757), .E(n6396), .CP(clk), .QN(n15517) );
  EDFD1 \Mem_reg[64][17]  ( .D(n24757), .E(n6395), .CP(clk), .QN(n5225) );
  EDFD1 \Mem_reg[63][17]  ( .D(n24757), .E(n6456), .CP(clk), .QN(n5177) );
  EDFD1 \Mem_reg[62][17]  ( .D(n24757), .E(n6455), .CP(clk), .QN(n5129) );
  EDFD1 \Mem_reg[61][17]  ( .D(n24757), .E(n6454), .CP(clk), .QN(n17978) );
  EDFD1 \Mem_reg[60][17]  ( .D(n24757), .E(n6453), .CP(clk), .QN(n17977) );
  EDFD1 \Mem_reg[59][17]  ( .D(n24757), .E(n6452), .CP(clk), .QN(n4985) );
  EDFD1 \Mem_reg[58][17]  ( .D(n24757), .E(n6451), .CP(clk), .QN(n4937) );
  EDFD1 \Mem_reg[57][17]  ( .D(n24757), .E(n6450), .CP(clk), .QN(n4889) );
  EDFD1 \Mem_reg[56][17]  ( .D(n24757), .E(n6449), .CP(clk), .QN(n4841) );
  EDFD1 \Mem_reg[55][17]  ( .D(n24757), .E(n6448), .CP(clk), .QN(n4793) );
  EDFD1 \Mem_reg[54][17]  ( .D(n24757), .E(n6447), .CP(clk), .QN(n15516) );
  EDFD1 \Mem_reg[53][17]  ( .D(n24757), .E(n6446), .CP(clk), .QN(n4697) );
  EDFD1 \Mem_reg[52][17]  ( .D(n24757), .E(n6445), .CP(clk), .Q(n27104) );
  EDFD1 \Mem_reg[51][17]  ( .D(n24757), .E(n6444), .CP(clk), .QN(n4601) );
  EDFD1 \Mem_reg[50][17]  ( .D(n24757), .E(n6443), .CP(clk), .QN(n4553) );
  EDFD1 \Mem_reg[49][17]  ( .D(n24757), .E(n6442), .CP(clk), .QN(n4505) );
  EDFD1 \Mem_reg[48][17]  ( .D(n24757), .E(n6441), .CP(clk), .QN(n4457) );
  EDFD1 \Mem_reg[47][17]  ( .D(n24757), .E(n6440), .CP(clk), .QN(n4409) );
  EDFD1 \Mem_reg[46][17]  ( .D(n24757), .E(n6439), .CP(clk), .QN(n4361) );
  EDFD1 \Mem_reg[43][17]  ( .D(n24757), .E(n6438), .CP(clk), .QN(n4313) );
  EDFD1 \Mem_reg[42][17]  ( .D(n24757), .E(n6437), .CP(clk), .QN(n4265) );
  EDFD1 \Mem_reg[41][17]  ( .D(n24757), .E(n6436), .CP(clk), .QN(n4217) );
  EDFD1 \Mem_reg[40][17]  ( .D(n24757), .E(n6435), .CP(clk), .QN(n4169) );
  EDFD1 \Mem_reg[39][17]  ( .D(n24757), .E(n6434), .CP(clk), .QN(n4121) );
  EDFD1 \Mem_reg[38][17]  ( .D(n24757), .E(n6433), .CP(clk), .QN(n4073) );
  EDFD1 \Mem_reg[37][17]  ( .D(n24757), .E(n6432), .CP(clk), .QN(n4025) );
  EDFD1 \Mem_reg[36][17]  ( .D(n24757), .E(n6431), .CP(clk), .QN(n3977) );
  EDFD1 \Mem_reg[35][17]  ( .D(n24757), .E(n6430), .CP(clk), .QN(n3929) );
  EDFD1 \Mem_reg[34][17]  ( .D(n24757), .E(n6429), .CP(clk), .QN(n3881) );
  EDFD1 \Mem_reg[33][17]  ( .D(n24757), .E(n6428), .CP(clk), .QN(n3833) );
  EDFD1 \Mem_reg[32][17]  ( .D(n24757), .E(n6427), .CP(clk), .QN(n3785) );
  EDFD1 \Mem_reg[31][17]  ( .D(n24757), .E(n6426), .CP(clk), .QN(n3737) );
  EDFD1 \Mem_reg[30][17]  ( .D(n24757), .E(n6425), .CP(clk), .QN(n3689) );
  EDFD1 \Mem_reg[29][17]  ( .D(n24757), .E(n6424), .CP(clk), .QN(n3641) );
  EDFD1 \Mem_reg[28][17]  ( .D(n24757), .E(n6423), .CP(clk), .QN(n3593) );
  EDFD1 \Mem_reg[27][17]  ( .D(n24757), .E(n6422), .CP(clk), .QN(n3545) );
  EDFD1 \Mem_reg[26][17]  ( .D(n24757), .E(n6421), .CP(clk), .QN(n3497) );
  EDFD1 \Mem_reg[25][17]  ( .D(n24757), .E(n6420), .CP(clk), .QN(n3449) );
  EDFD1 \Mem_reg[24][17]  ( .D(n24757), .E(n6463), .CP(clk), .QN(n3401) );
  EDFD1 \Mem_reg[23][17]  ( .D(n24757), .E(n6464), .CP(clk), .QN(n3353) );
  EDFD1 \Mem_reg[22][17]  ( .D(n24757), .E(n6465), .CP(clk), .QN(n3305) );
  EDFD1 \Mem_reg[21][17]  ( .D(n24757), .E(n6466), .CP(clk), .QN(n3257) );
  EDFD1 \Mem_reg[20][17]  ( .D(n24757), .E(n6467), .CP(clk), .QN(n3209) );
  EDFD1 \Mem_reg[19][17]  ( .D(n24757), .E(n6468), .CP(clk), .QN(n3161) );
  EDFD1 \Mem_reg[18][17]  ( .D(n24757), .E(n6469), .CP(clk), .QN(n3113) );
  EDFD1 \Mem_reg[17][17]  ( .D(n24757), .E(n6470), .CP(clk), .QN(n3065) );
  EDFD1 \Mem_reg[16][17]  ( .D(n24757), .E(n6471), .CP(clk), .QN(n3017) );
  EDFD1 \Mem_reg[15][17]  ( .D(n24757), .E(n6472), .CP(clk), .QN(n2969) );
  EDFD1 \Mem_reg[14][17]  ( .D(n24757), .E(n24720), .CP(clk), .QN(n2921) );
  EDFD1 \Mem_reg[13][17]  ( .D(n24757), .E(n24709), .CP(clk), .QN(n2873) );
  EDFD1 \Mem_reg[12][17]  ( .D(n24757), .E(n24717), .CP(clk), .QN(n2825) );
  EDFD1 \Mem_reg[11][17]  ( .D(n24757), .E(n24707), .CP(clk), .QN(n2777) );
  EDFD1 \Mem_reg[10][17]  ( .D(n24757), .E(n6477), .CP(clk), .QN(n2729) );
  EDFD1 \Mem_reg[9][17]  ( .D(n24757), .E(n24708), .CP(clk), .QN(n2681) );
  EDFD1 \Mem_reg[8][17]  ( .D(n24757), .E(n15642), .CP(clk), .QN(n2633) );
  EDFD1 \Mem_reg[7][17]  ( .D(n24757), .E(n24718), .CP(clk), .QN(n2585) );
  EDFD1 \Mem_reg[6][17]  ( .D(n24757), .E(n24716), .CP(clk), .QN(n2537) );
  EDFD1 \Mem_reg[5][17]  ( .D(n24757), .E(n24719), .CP(clk), .QN(n2489) );
  EDFD1 \Mem_reg[4][17]  ( .D(n24757), .E(n24706), .CP(clk), .QN(n2441) );
  EDFD1 \Mem_reg[3][17]  ( .D(n24757), .E(n24721), .CP(clk), .QN(n2393) );
  EDFD1 \Mem_reg[2][17]  ( .D(n24757), .E(n6460), .CP(clk), .QN(n2345) );
  EDFD1 \Mem_reg[1][17]  ( .D(n24757), .E(n24703), .CP(clk), .QN(n2297) );
  EDFD1 \Mem_reg[0][17]  ( .D(n24757), .E(n24705), .CP(clk), .QN(n2249) );
  EDFD1 \Mem_reg[88][16]  ( .D(n24755), .E(n6419), .CP(clk), .Q(n27101) );
  EDFD1 \Mem_reg[87][16]  ( .D(n24755), .E(n6418), .CP(clk), .QN(n6330) );
  EDFD1 \Mem_reg[86][16]  ( .D(n24755), .E(n6417), .CP(clk), .QN(n24607) );
  EDFD1 \Mem_reg[85][16]  ( .D(n24755), .E(n6416), .CP(clk), .QN(n6234) );
  EDFD1 \Mem_reg[84][16]  ( .D(n24755), .E(n6415), .CP(clk), .QN(n6186) );
  EDFD1 \Mem_reg[83][16]  ( .D(n24755), .E(n6414), .CP(clk), .QN(n6138) );
  EDFD1 \Mem_reg[82][16]  ( .D(n24755), .E(n6413), .CP(clk), .QN(n6090) );
  EDFD1 \Mem_reg[81][16]  ( .D(n24755), .E(n6412), .CP(clk), .QN(n6042) );
  EDFD1 \Mem_reg[80][16]  ( .D(n24755), .E(n6411), .CP(clk), .QN(n5994) );
  EDFD1 \Mem_reg[79][16]  ( .D(n24755), .E(n6410), .CP(clk), .QN(n5946) );
  EDFD1 \Mem_reg[78][16]  ( .D(n24755), .E(n6409), .CP(clk), .QN(n5898) );
  EDFD1 \Mem_reg[77][16]  ( .D(n24755), .E(n6408), .CP(clk), .QN(n5850) );
  EDFD1 \Mem_reg[76][16]  ( .D(n24755), .E(n6407), .CP(clk), .QN(n5802) );
  EDFD1 \Mem_reg[75][16]  ( .D(n24755), .E(n6406), .CP(clk), .QN(n27102) );
  EDFD1 \Mem_reg[74][16]  ( .D(n24755), .E(n6405), .CP(clk), .QN(n5706) );
  EDFD1 \Mem_reg[73][16]  ( .D(n24755), .E(n6404), .CP(clk), .QN(n27103) );
  EDFD1 \Mem_reg[72][16]  ( .D(n24755), .E(n6403), .CP(clk), .QN(n5610) );
  EDFD1 \Mem_reg[71][16]  ( .D(n24755), .E(n6402), .CP(clk), .QN(n5562) );
  EDFD1 \Mem_reg[70][16]  ( .D(n24755), .E(n6401), .CP(clk), .QN(n5514) );
  EDFD1 \Mem_reg[69][16]  ( .D(n24755), .E(n6400), .CP(clk), .QN(n5466) );
  EDFD1 \Mem_reg[68][16]  ( .D(n24755), .E(n6399), .CP(clk), .QN(n5418) );
  EDFD1 \Mem_reg[67][16]  ( .D(n24755), .E(n6398), .CP(clk), .QN(n5370) );
  EDFD1 \Mem_reg[66][16]  ( .D(n24755), .E(n6397), .CP(clk), .QN(n5322) );
  EDFD1 \Mem_reg[65][16]  ( .D(n24755), .E(n6396), .CP(clk), .QN(n15513) );
  EDFD1 \Mem_reg[64][16]  ( .D(n24755), .E(n6395), .CP(clk), .QN(n5226) );
  EDFD1 \Mem_reg[63][16]  ( .D(n24755), .E(n6456), .CP(clk), .QN(n5178) );
  EDFD1 \Mem_reg[62][16]  ( .D(n24755), .E(n6455), .CP(clk), .QN(n5130) );
  EDFD1 \Mem_reg[61][16]  ( .D(n24755), .E(n6454), .CP(clk), .QN(n17975) );
  EDFD1 \Mem_reg[60][16]  ( .D(n24755), .E(n6453), .CP(clk), .QN(n17974) );
  EDFD1 \Mem_reg[59][16]  ( .D(n24755), .E(n6452), .CP(clk), .QN(n4986) );
  EDFD1 \Mem_reg[58][16]  ( .D(n24755), .E(n6451), .CP(clk), .QN(n4938) );
  EDFD1 \Mem_reg[57][16]  ( .D(n24755), .E(n6450), .CP(clk), .QN(n4890) );
  EDFD1 \Mem_reg[56][16]  ( .D(n24755), .E(n6449), .CP(clk), .QN(n4842) );
  EDFD1 \Mem_reg[55][16]  ( .D(n24755), .E(n6448), .CP(clk), .QN(n4794) );
  EDFD1 \Mem_reg[54][16]  ( .D(n24755), .E(n6447), .CP(clk), .QN(n15512) );
  EDFD1 \Mem_reg[53][16]  ( .D(n24755), .E(n6446), .CP(clk), .QN(n4698) );
  EDFD1 \Mem_reg[52][16]  ( .D(n24755), .E(n6445), .CP(clk), .Q(n27100) );
  EDFD1 \Mem_reg[51][16]  ( .D(n24755), .E(n6444), .CP(clk), .QN(n4602) );
  EDFD1 \Mem_reg[50][16]  ( .D(n24755), .E(n6443), .CP(clk), .QN(n4554) );
  EDFD1 \Mem_reg[49][16]  ( .D(n24755), .E(n6442), .CP(clk), .QN(n4506) );
  EDFD1 \Mem_reg[48][16]  ( .D(n24755), .E(n6441), .CP(clk), .QN(n4458) );
  EDFD1 \Mem_reg[47][16]  ( .D(n24755), .E(n6440), .CP(clk), .QN(n4410) );
  EDFD1 \Mem_reg[46][16]  ( .D(n24755), .E(n6439), .CP(clk), .QN(n4362) );
  EDFD1 \Mem_reg[43][16]  ( .D(n24755), .E(n6438), .CP(clk), .QN(n4314) );
  EDFD1 \Mem_reg[42][16]  ( .D(n24755), .E(n6437), .CP(clk), .QN(n4266) );
  EDFD1 \Mem_reg[41][16]  ( .D(n24755), .E(n6436), .CP(clk), .QN(n4218) );
  EDFD1 \Mem_reg[40][16]  ( .D(n24755), .E(n6435), .CP(clk), .QN(n4170) );
  EDFD1 \Mem_reg[39][16]  ( .D(n24755), .E(n6434), .CP(clk), .QN(n4122) );
  EDFD1 \Mem_reg[38][16]  ( .D(n24755), .E(n6433), .CP(clk), .QN(n4074) );
  EDFD1 \Mem_reg[37][16]  ( .D(n24755), .E(n6432), .CP(clk), .QN(n4026) );
  EDFD1 \Mem_reg[36][16]  ( .D(n24755), .E(n6431), .CP(clk), .QN(n3978) );
  EDFD1 \Mem_reg[35][16]  ( .D(n24755), .E(n6430), .CP(clk), .QN(n3930) );
  EDFD1 \Mem_reg[34][16]  ( .D(n24755), .E(n6429), .CP(clk), .QN(n3882) );
  EDFD1 \Mem_reg[33][16]  ( .D(n24755), .E(n6428), .CP(clk), .QN(n3834) );
  EDFD1 \Mem_reg[32][16]  ( .D(n24755), .E(n6427), .CP(clk), .QN(n3786) );
  EDFD1 \Mem_reg[31][16]  ( .D(n24755), .E(n6426), .CP(clk), .QN(n3738) );
  EDFD1 \Mem_reg[30][16]  ( .D(n24755), .E(n6425), .CP(clk), .QN(n3690) );
  EDFD1 \Mem_reg[29][16]  ( .D(n24755), .E(n6424), .CP(clk), .QN(n3642) );
  EDFD1 \Mem_reg[28][16]  ( .D(n24755), .E(n6423), .CP(clk), .QN(n3594) );
  EDFD1 \Mem_reg[27][16]  ( .D(n24755), .E(n6422), .CP(clk), .QN(n3546) );
  EDFD1 \Mem_reg[26][16]  ( .D(n24755), .E(n6421), .CP(clk), .QN(n3498) );
  EDFD1 \Mem_reg[25][16]  ( .D(n24755), .E(n6420), .CP(clk), .QN(n3450) );
  EDFD1 \Mem_reg[24][16]  ( .D(n24755), .E(n6463), .CP(clk), .QN(n3402) );
  EDFD1 \Mem_reg[23][16]  ( .D(n24755), .E(n6464), .CP(clk), .QN(n3354) );
  EDFD1 \Mem_reg[22][16]  ( .D(n24755), .E(n6465), .CP(clk), .QN(n3306) );
  EDFD1 \Mem_reg[21][16]  ( .D(n24755), .E(n6466), .CP(clk), .QN(n3258) );
  EDFD1 \Mem_reg[20][16]  ( .D(n24755), .E(n6467), .CP(clk), .QN(n3210) );
  EDFD1 \Mem_reg[19][16]  ( .D(n24755), .E(n6468), .CP(clk), .QN(n3162) );
  EDFD1 \Mem_reg[18][16]  ( .D(n24755), .E(n6469), .CP(clk), .QN(n3114) );
  EDFD1 \Mem_reg[17][16]  ( .D(n24755), .E(n6470), .CP(clk), .QN(n3066) );
  EDFD1 \Mem_reg[16][16]  ( .D(n24755), .E(n6471), .CP(clk), .QN(n3018) );
  EDFD1 \Mem_reg[15][16]  ( .D(n24755), .E(n6472), .CP(clk), .QN(n2970) );
  EDFD1 \Mem_reg[14][16]  ( .D(n24755), .E(n24720), .CP(clk), .QN(n2922) );
  EDFD1 \Mem_reg[13][16]  ( .D(n24755), .E(n24709), .CP(clk), .QN(n2874) );
  EDFD1 \Mem_reg[12][16]  ( .D(n24755), .E(n24717), .CP(clk), .QN(n2826) );
  EDFD1 \Mem_reg[11][16]  ( .D(n24755), .E(n24707), .CP(clk), .QN(n2778) );
  EDFD1 \Mem_reg[10][16]  ( .D(n24755), .E(n6477), .CP(clk), .QN(n2730) );
  EDFD1 \Mem_reg[9][16]  ( .D(n24755), .E(n24708), .CP(clk), .QN(n2682) );
  EDFD1 \Mem_reg[8][16]  ( .D(n24755), .E(n15642), .CP(clk), .QN(n2634) );
  EDFD1 \Mem_reg[7][16]  ( .D(n24755), .E(n24718), .CP(clk), .QN(n2586) );
  EDFD1 \Mem_reg[6][16]  ( .D(n24755), .E(n24716), .CP(clk), .QN(n2538) );
  EDFD1 \Mem_reg[5][16]  ( .D(n24755), .E(n24719), .CP(clk), .QN(n2490) );
  EDFD1 \Mem_reg[4][16]  ( .D(n24755), .E(n24706), .CP(clk), .QN(n2442) );
  EDFD1 \Mem_reg[3][16]  ( .D(n24755), .E(n24721), .CP(clk), .QN(n2394) );
  EDFD1 \Mem_reg[2][16]  ( .D(n24755), .E(n6460), .CP(clk), .QN(n2346) );
  EDFD1 \Mem_reg[1][16]  ( .D(n24755), .E(n24703), .CP(clk), .QN(n2298) );
  EDFD1 \Mem_reg[0][16]  ( .D(n24755), .E(n24705), .CP(clk), .QN(n2250) );
  EDFD1 \Mem_reg[88][15]  ( .D(n24753), .E(n6419), .CP(clk), .Q(n27097) );
  EDFD1 \Mem_reg[87][15]  ( .D(n24753), .E(n6418), .CP(clk), .QN(n6331) );
  EDFD1 \Mem_reg[86][15]  ( .D(n24753), .E(n6417), .CP(clk), .QN(n24604) );
  EDFD1 \Mem_reg[85][15]  ( .D(n24753), .E(n6416), .CP(clk), .QN(n6235) );
  EDFD1 \Mem_reg[84][15]  ( .D(n24753), .E(n6415), .CP(clk), .QN(n6187) );
  EDFD1 \Mem_reg[83][15]  ( .D(n24753), .E(n6414), .CP(clk), .QN(n6139) );
  EDFD1 \Mem_reg[82][15]  ( .D(n24753), .E(n6413), .CP(clk), .QN(n6091) );
  EDFD1 \Mem_reg[81][15]  ( .D(n24753), .E(n6412), .CP(clk), .QN(n6043) );
  EDFD1 \Mem_reg[80][15]  ( .D(n24753), .E(n6411), .CP(clk), .QN(n5995) );
  EDFD1 \Mem_reg[79][15]  ( .D(n24753), .E(n6410), .CP(clk), .QN(n5947) );
  EDFD1 \Mem_reg[78][15]  ( .D(n24753), .E(n6409), .CP(clk), .QN(n5899) );
  EDFD1 \Mem_reg[77][15]  ( .D(n24753), .E(n6408), .CP(clk), .QN(n5851) );
  EDFD1 \Mem_reg[76][15]  ( .D(n24753), .E(n6407), .CP(clk), .QN(n5803) );
  EDFD1 \Mem_reg[75][15]  ( .D(n24753), .E(n6406), .CP(clk), .QN(n27098) );
  EDFD1 \Mem_reg[74][15]  ( .D(n24753), .E(n6405), .CP(clk), .QN(n5707) );
  EDFD1 \Mem_reg[73][15]  ( .D(n24753), .E(n6404), .CP(clk), .QN(n27099) );
  EDFD1 \Mem_reg[72][15]  ( .D(n24753), .E(n6403), .CP(clk), .QN(n5611) );
  EDFD1 \Mem_reg[71][15]  ( .D(n24753), .E(n6402), .CP(clk), .QN(n5563) );
  EDFD1 \Mem_reg[70][15]  ( .D(n24753), .E(n6401), .CP(clk), .QN(n5515) );
  EDFD1 \Mem_reg[69][15]  ( .D(n24753), .E(n6400), .CP(clk), .QN(n5467) );
  EDFD1 \Mem_reg[68][15]  ( .D(n24753), .E(n6399), .CP(clk), .QN(n5419) );
  EDFD1 \Mem_reg[67][15]  ( .D(n24753), .E(n6398), .CP(clk), .QN(n5371) );
  EDFD1 \Mem_reg[66][15]  ( .D(n24753), .E(n6397), .CP(clk), .QN(n5323) );
  EDFD1 \Mem_reg[65][15]  ( .D(n24753), .E(n6396), .CP(clk), .QN(n15509) );
  EDFD1 \Mem_reg[64][15]  ( .D(n24753), .E(n6395), .CP(clk), .QN(n5227) );
  EDFD1 \Mem_reg[63][15]  ( .D(n24753), .E(n6456), .CP(clk), .QN(n5179) );
  EDFD1 \Mem_reg[62][15]  ( .D(n24753), .E(n6455), .CP(clk), .QN(n5131) );
  EDFD1 \Mem_reg[61][15]  ( .D(n24753), .E(n6454), .CP(clk), .QN(n17972) );
  EDFD1 \Mem_reg[60][15]  ( .D(n24753), .E(n6453), .CP(clk), .QN(n17971) );
  EDFD1 \Mem_reg[59][15]  ( .D(n24753), .E(n6452), .CP(clk), .QN(n4987) );
  EDFD1 \Mem_reg[58][15]  ( .D(n24753), .E(n6451), .CP(clk), .QN(n4939) );
  EDFD1 \Mem_reg[57][15]  ( .D(n24753), .E(n6450), .CP(clk), .QN(n4891) );
  EDFD1 \Mem_reg[56][15]  ( .D(n24753), .E(n6449), .CP(clk), .QN(n4843) );
  EDFD1 \Mem_reg[55][15]  ( .D(n24753), .E(n6448), .CP(clk), .QN(n4795) );
  EDFD1 \Mem_reg[54][15]  ( .D(n24753), .E(n6447), .CP(clk), .QN(n15508) );
  EDFD1 \Mem_reg[53][15]  ( .D(n24753), .E(n6446), .CP(clk), .QN(n4699) );
  EDFD1 \Mem_reg[52][15]  ( .D(n24753), .E(n6445), .CP(clk), .Q(n27096) );
  EDFD1 \Mem_reg[51][15]  ( .D(n24753), .E(n6444), .CP(clk), .QN(n4603) );
  EDFD1 \Mem_reg[50][15]  ( .D(n24753), .E(n6443), .CP(clk), .QN(n4555) );
  EDFD1 \Mem_reg[49][15]  ( .D(n24753), .E(n6442), .CP(clk), .QN(n4507) );
  EDFD1 \Mem_reg[48][15]  ( .D(n24753), .E(n6441), .CP(clk), .QN(n4459) );
  EDFD1 \Mem_reg[47][15]  ( .D(n24753), .E(n6440), .CP(clk), .QN(n4411) );
  EDFD1 \Mem_reg[46][15]  ( .D(n24753), .E(n6439), .CP(clk), .QN(n4363) );
  EDFD1 \Mem_reg[43][15]  ( .D(n24753), .E(n6438), .CP(clk), .QN(n4315) );
  EDFD1 \Mem_reg[42][15]  ( .D(n24753), .E(n6437), .CP(clk), .QN(n4267) );
  EDFD1 \Mem_reg[41][15]  ( .D(n24753), .E(n6436), .CP(clk), .QN(n4219) );
  EDFD1 \Mem_reg[40][15]  ( .D(n24753), .E(n6435), .CP(clk), .QN(n4171) );
  EDFD1 \Mem_reg[39][15]  ( .D(n24753), .E(n6434), .CP(clk), .QN(n4123) );
  EDFD1 \Mem_reg[38][15]  ( .D(n24753), .E(n6433), .CP(clk), .QN(n4075) );
  EDFD1 \Mem_reg[37][15]  ( .D(n24753), .E(n6432), .CP(clk), .QN(n4027) );
  EDFD1 \Mem_reg[36][15]  ( .D(n24753), .E(n6431), .CP(clk), .QN(n3979) );
  EDFD1 \Mem_reg[35][15]  ( .D(n24753), .E(n6430), .CP(clk), .QN(n3931) );
  EDFD1 \Mem_reg[34][15]  ( .D(n24753), .E(n6429), .CP(clk), .QN(n3883) );
  EDFD1 \Mem_reg[33][15]  ( .D(n24753), .E(n6428), .CP(clk), .QN(n3835) );
  EDFD1 \Mem_reg[32][15]  ( .D(n24753), .E(n6427), .CP(clk), .QN(n3787) );
  EDFD1 \Mem_reg[31][15]  ( .D(n24753), .E(n6426), .CP(clk), .QN(n3739) );
  EDFD1 \Mem_reg[30][15]  ( .D(n24753), .E(n6425), .CP(clk), .QN(n3691) );
  EDFD1 \Mem_reg[29][15]  ( .D(n24753), .E(n6424), .CP(clk), .QN(n3643) );
  EDFD1 \Mem_reg[28][15]  ( .D(n24753), .E(n6423), .CP(clk), .QN(n3595) );
  EDFD1 \Mem_reg[27][15]  ( .D(n24753), .E(n6422), .CP(clk), .QN(n3547) );
  EDFD1 \Mem_reg[26][15]  ( .D(n24753), .E(n6421), .CP(clk), .QN(n3499) );
  EDFD1 \Mem_reg[25][15]  ( .D(n24753), .E(n6420), .CP(clk), .QN(n3451) );
  EDFD1 \Mem_reg[24][15]  ( .D(n24753), .E(n6463), .CP(clk), .QN(n3403) );
  EDFD1 \Mem_reg[23][15]  ( .D(n24753), .E(n6464), .CP(clk), .QN(n3355) );
  EDFD1 \Mem_reg[22][15]  ( .D(n24753), .E(n6465), .CP(clk), .QN(n3307) );
  EDFD1 \Mem_reg[21][15]  ( .D(n24753), .E(n6466), .CP(clk), .QN(n3259) );
  EDFD1 \Mem_reg[20][15]  ( .D(n24753), .E(n6467), .CP(clk), .QN(n3211) );
  EDFD1 \Mem_reg[19][15]  ( .D(n24753), .E(n6468), .CP(clk), .QN(n3163) );
  EDFD1 \Mem_reg[18][15]  ( .D(n24753), .E(n6469), .CP(clk), .QN(n3115) );
  EDFD1 \Mem_reg[17][15]  ( .D(n24753), .E(n6470), .CP(clk), .QN(n3067) );
  EDFD1 \Mem_reg[16][15]  ( .D(n24753), .E(n6471), .CP(clk), .QN(n3019) );
  EDFD1 \Mem_reg[15][15]  ( .D(n24753), .E(n6472), .CP(clk), .QN(n2971) );
  EDFD1 \Mem_reg[14][15]  ( .D(n24753), .E(n24720), .CP(clk), .QN(n2923) );
  EDFD1 \Mem_reg[13][15]  ( .D(n24753), .E(n24709), .CP(clk), .QN(n2875) );
  EDFD1 \Mem_reg[12][15]  ( .D(n24753), .E(n24717), .CP(clk), .QN(n2827) );
  EDFD1 \Mem_reg[11][15]  ( .D(n24753), .E(n24707), .CP(clk), .QN(n2779) );
  EDFD1 \Mem_reg[10][15]  ( .D(n24753), .E(n6477), .CP(clk), .QN(n2731) );
  EDFD1 \Mem_reg[9][15]  ( .D(n24753), .E(n24708), .CP(clk), .QN(n2683) );
  EDFD1 \Mem_reg[8][15]  ( .D(n24753), .E(n15642), .CP(clk), .QN(n2635) );
  EDFD1 \Mem_reg[7][15]  ( .D(n24753), .E(n24718), .CP(clk), .QN(n2587) );
  EDFD1 \Mem_reg[6][15]  ( .D(n24753), .E(n24716), .CP(clk), .QN(n2539) );
  EDFD1 \Mem_reg[5][15]  ( .D(n24753), .E(n24719), .CP(clk), .QN(n2491) );
  EDFD1 \Mem_reg[4][15]  ( .D(n24753), .E(n24706), .CP(clk), .QN(n2443) );
  EDFD1 \Mem_reg[3][15]  ( .D(n24753), .E(n24721), .CP(clk), .QN(n2395) );
  EDFD1 \Mem_reg[2][15]  ( .D(n24753), .E(n6460), .CP(clk), .QN(n2347) );
  EDFD1 \Mem_reg[1][15]  ( .D(n24753), .E(n24703), .CP(clk), .QN(n2299) );
  EDFD1 \Mem_reg[0][15]  ( .D(n24753), .E(n24705), .CP(clk), .QN(n2251) );
  EDFD1 \Mem_reg[88][14]  ( .D(n24751), .E(n6419), .CP(clk), .Q(n27093) );
  EDFD1 \Mem_reg[87][14]  ( .D(n24751), .E(n6418), .CP(clk), .QN(n6332) );
  EDFD1 \Mem_reg[86][14]  ( .D(n24751), .E(n6417), .CP(clk), .QN(n24601) );
  EDFD1 \Mem_reg[85][14]  ( .D(n24751), .E(n6416), .CP(clk), .QN(n6236) );
  EDFD1 \Mem_reg[84][14]  ( .D(n24751), .E(n6415), .CP(clk), .QN(n6188) );
  EDFD1 \Mem_reg[83][14]  ( .D(n24751), .E(n6414), .CP(clk), .QN(n6140) );
  EDFD1 \Mem_reg[82][14]  ( .D(n24751), .E(n6413), .CP(clk), .QN(n6092) );
  EDFD1 \Mem_reg[81][14]  ( .D(n24751), .E(n6412), .CP(clk), .QN(n6044) );
  EDFD1 \Mem_reg[80][14]  ( .D(n24751), .E(n6411), .CP(clk), .QN(n5996) );
  EDFD1 \Mem_reg[79][14]  ( .D(n24751), .E(n6410), .CP(clk), .QN(n5948) );
  EDFD1 \Mem_reg[78][14]  ( .D(n24751), .E(n6409), .CP(clk), .QN(n5900) );
  EDFD1 \Mem_reg[77][14]  ( .D(n24751), .E(n6408), .CP(clk), .QN(n5852) );
  EDFD1 \Mem_reg[76][14]  ( .D(n24751), .E(n6407), .CP(clk), .QN(n5804) );
  EDFD1 \Mem_reg[75][14]  ( .D(n24751), .E(n6406), .CP(clk), .QN(n27094) );
  EDFD1 \Mem_reg[74][14]  ( .D(n24751), .E(n6405), .CP(clk), .QN(n5708) );
  EDFD1 \Mem_reg[73][14]  ( .D(n24751), .E(n6404), .CP(clk), .QN(n27095) );
  EDFD1 \Mem_reg[72][14]  ( .D(n24751), .E(n6403), .CP(clk), .QN(n5612) );
  EDFD1 \Mem_reg[71][14]  ( .D(n24751), .E(n6402), .CP(clk), .QN(n5564) );
  EDFD1 \Mem_reg[70][14]  ( .D(n24751), .E(n6401), .CP(clk), .QN(n5516) );
  EDFD1 \Mem_reg[69][14]  ( .D(n24751), .E(n6400), .CP(clk), .QN(n5468) );
  EDFD1 \Mem_reg[68][14]  ( .D(n24751), .E(n6399), .CP(clk), .QN(n5420) );
  EDFD1 \Mem_reg[67][14]  ( .D(n24751), .E(n6398), .CP(clk), .QN(n5372) );
  EDFD1 \Mem_reg[66][14]  ( .D(n24751), .E(n6397), .CP(clk), .QN(n5324) );
  EDFD1 \Mem_reg[65][14]  ( .D(n24751), .E(n6396), .CP(clk), .QN(n15505) );
  EDFD1 \Mem_reg[64][14]  ( .D(n24751), .E(n6395), .CP(clk), .QN(n5228) );
  EDFD1 \Mem_reg[63][14]  ( .D(n24751), .E(n6456), .CP(clk), .QN(n5180) );
  EDFD1 \Mem_reg[62][14]  ( .D(n24751), .E(n6455), .CP(clk), .QN(n5132) );
  EDFD1 \Mem_reg[61][14]  ( .D(n24751), .E(n6454), .CP(clk), .QN(n17969) );
  EDFD1 \Mem_reg[60][14]  ( .D(n24751), .E(n6453), .CP(clk), .QN(n17968) );
  EDFD1 \Mem_reg[59][14]  ( .D(n24751), .E(n6452), .CP(clk), .QN(n4988) );
  EDFD1 \Mem_reg[58][14]  ( .D(n24751), .E(n6451), .CP(clk), .QN(n4940) );
  EDFD1 \Mem_reg[57][14]  ( .D(n24751), .E(n6450), .CP(clk), .QN(n4892) );
  EDFD1 \Mem_reg[56][14]  ( .D(n24751), .E(n6449), .CP(clk), .QN(n4844) );
  EDFD1 \Mem_reg[55][14]  ( .D(n24751), .E(n6448), .CP(clk), .QN(n4796) );
  EDFD1 \Mem_reg[54][14]  ( .D(n24751), .E(n6447), .CP(clk), .QN(n15504) );
  EDFD1 \Mem_reg[53][14]  ( .D(n24751), .E(n6446), .CP(clk), .QN(n4700) );
  EDFD1 \Mem_reg[52][14]  ( .D(n24751), .E(n6445), .CP(clk), .Q(n27092) );
  EDFD1 \Mem_reg[51][14]  ( .D(n24751), .E(n6444), .CP(clk), .QN(n4604) );
  EDFD1 \Mem_reg[50][14]  ( .D(n24751), .E(n6443), .CP(clk), .QN(n4556) );
  EDFD1 \Mem_reg[49][14]  ( .D(n24751), .E(n6442), .CP(clk), .QN(n4508) );
  EDFD1 \Mem_reg[48][14]  ( .D(n24751), .E(n6441), .CP(clk), .QN(n4460) );
  EDFD1 \Mem_reg[47][14]  ( .D(n24751), .E(n6440), .CP(clk), .QN(n4412) );
  EDFD1 \Mem_reg[46][14]  ( .D(n24751), .E(n6439), .CP(clk), .QN(n4364) );
  EDFD1 \Mem_reg[43][14]  ( .D(n24751), .E(n6438), .CP(clk), .QN(n4316) );
  EDFD1 \Mem_reg[42][14]  ( .D(n24751), .E(n6437), .CP(clk), .QN(n4268) );
  EDFD1 \Mem_reg[41][14]  ( .D(n24751), .E(n6436), .CP(clk), .QN(n4220) );
  EDFD1 \Mem_reg[40][14]  ( .D(n24751), .E(n6435), .CP(clk), .QN(n4172) );
  EDFD1 \Mem_reg[39][14]  ( .D(n24751), .E(n6434), .CP(clk), .QN(n4124) );
  EDFD1 \Mem_reg[38][14]  ( .D(n24751), .E(n6433), .CP(clk), .QN(n4076) );
  EDFD1 \Mem_reg[37][14]  ( .D(n24751), .E(n6432), .CP(clk), .QN(n4028) );
  EDFD1 \Mem_reg[36][14]  ( .D(n24751), .E(n6431), .CP(clk), .QN(n3980) );
  EDFD1 \Mem_reg[35][14]  ( .D(n24751), .E(n6430), .CP(clk), .QN(n3932) );
  EDFD1 \Mem_reg[34][14]  ( .D(n24751), .E(n6429), .CP(clk), .QN(n3884) );
  EDFD1 \Mem_reg[33][14]  ( .D(n24751), .E(n6428), .CP(clk), .QN(n3836) );
  EDFD1 \Mem_reg[32][14]  ( .D(n24751), .E(n6427), .CP(clk), .QN(n3788) );
  EDFD1 \Mem_reg[31][14]  ( .D(n24751), .E(n6426), .CP(clk), .QN(n3740) );
  EDFD1 \Mem_reg[30][14]  ( .D(n24751), .E(n6425), .CP(clk), .QN(n3692) );
  EDFD1 \Mem_reg[29][14]  ( .D(n24751), .E(n6424), .CP(clk), .QN(n3644) );
  EDFD1 \Mem_reg[28][14]  ( .D(n24751), .E(n6423), .CP(clk), .QN(n3596) );
  EDFD1 \Mem_reg[27][14]  ( .D(n24751), .E(n6422), .CP(clk), .QN(n3548) );
  EDFD1 \Mem_reg[26][14]  ( .D(n24751), .E(n6421), .CP(clk), .QN(n3500) );
  EDFD1 \Mem_reg[25][14]  ( .D(n24751), .E(n6420), .CP(clk), .QN(n3452) );
  EDFD1 \Mem_reg[24][14]  ( .D(n24751), .E(n6463), .CP(clk), .QN(n3404) );
  EDFD1 \Mem_reg[23][14]  ( .D(n24751), .E(n6464), .CP(clk), .QN(n3356) );
  EDFD1 \Mem_reg[22][14]  ( .D(n24751), .E(n6465), .CP(clk), .QN(n3308) );
  EDFD1 \Mem_reg[21][14]  ( .D(n24751), .E(n6466), .CP(clk), .QN(n3260) );
  EDFD1 \Mem_reg[20][14]  ( .D(n24751), .E(n6467), .CP(clk), .QN(n3212) );
  EDFD1 \Mem_reg[19][14]  ( .D(n24751), .E(n6468), .CP(clk), .QN(n3164) );
  EDFD1 \Mem_reg[18][14]  ( .D(n24751), .E(n6469), .CP(clk), .QN(n3116) );
  EDFD1 \Mem_reg[17][14]  ( .D(n24751), .E(n6470), .CP(clk), .QN(n3068) );
  EDFD1 \Mem_reg[16][14]  ( .D(n24751), .E(n6471), .CP(clk), .QN(n3020) );
  EDFD1 \Mem_reg[15][14]  ( .D(n24751), .E(n6472), .CP(clk), .QN(n2972) );
  EDFD1 \Mem_reg[14][14]  ( .D(n24751), .E(n24720), .CP(clk), .QN(n2924) );
  EDFD1 \Mem_reg[13][14]  ( .D(n24751), .E(n24709), .CP(clk), .QN(n2876) );
  EDFD1 \Mem_reg[12][14]  ( .D(n24751), .E(n24717), .CP(clk), .QN(n2828) );
  EDFD1 \Mem_reg[11][14]  ( .D(n24751), .E(n24707), .CP(clk), .QN(n2780) );
  EDFD1 \Mem_reg[10][14]  ( .D(n24751), .E(n6477), .CP(clk), .QN(n2732) );
  EDFD1 \Mem_reg[9][14]  ( .D(n24751), .E(n24708), .CP(clk), .QN(n2684) );
  EDFD1 \Mem_reg[8][14]  ( .D(n24751), .E(n15642), .CP(clk), .QN(n2636) );
  EDFD1 \Mem_reg[7][14]  ( .D(n24751), .E(n24718), .CP(clk), .QN(n2588) );
  EDFD1 \Mem_reg[6][14]  ( .D(n24751), .E(n24716), .CP(clk), .QN(n2540) );
  EDFD1 \Mem_reg[5][14]  ( .D(n24751), .E(n24719), .CP(clk), .QN(n2492) );
  EDFD1 \Mem_reg[4][14]  ( .D(n24751), .E(n24706), .CP(clk), .QN(n2444) );
  EDFD1 \Mem_reg[3][14]  ( .D(n24751), .E(n24721), .CP(clk), .QN(n2396) );
  EDFD1 \Mem_reg[2][14]  ( .D(n24751), .E(n6460), .CP(clk), .QN(n2348) );
  EDFD1 \Mem_reg[1][14]  ( .D(n24751), .E(n24703), .CP(clk), .QN(n2300) );
  EDFD1 \Mem_reg[0][14]  ( .D(n24751), .E(n24705), .CP(clk), .QN(n2252) );
  EDFD1 \Mem_reg[88][13]  ( .D(n24749), .E(n6419), .CP(clk), .Q(n27089) );
  EDFD1 \Mem_reg[87][13]  ( .D(n24749), .E(n6418), .CP(clk), .QN(n6333) );
  EDFD1 \Mem_reg[86][13]  ( .D(n24749), .E(n6417), .CP(clk), .QN(n24598) );
  EDFD1 \Mem_reg[85][13]  ( .D(n24749), .E(n6416), .CP(clk), .QN(n6237) );
  EDFD1 \Mem_reg[84][13]  ( .D(n24749), .E(n6415), .CP(clk), .QN(n6189) );
  EDFD1 \Mem_reg[83][13]  ( .D(n24749), .E(n6414), .CP(clk), .QN(n6141) );
  EDFD1 \Mem_reg[82][13]  ( .D(n24749), .E(n6413), .CP(clk), .QN(n6093) );
  EDFD1 \Mem_reg[81][13]  ( .D(n24749), .E(n6412), .CP(clk), .QN(n6045) );
  EDFD1 \Mem_reg[80][13]  ( .D(n24749), .E(n6411), .CP(clk), .QN(n5997) );
  EDFD1 \Mem_reg[79][13]  ( .D(n24749), .E(n6410), .CP(clk), .QN(n5949) );
  EDFD1 \Mem_reg[78][13]  ( .D(n24749), .E(n6409), .CP(clk), .QN(n5901) );
  EDFD1 \Mem_reg[77][13]  ( .D(n24749), .E(n6408), .CP(clk), .QN(n5853) );
  EDFD1 \Mem_reg[76][13]  ( .D(n24749), .E(n6407), .CP(clk), .QN(n5805) );
  EDFD1 \Mem_reg[75][13]  ( .D(n24749), .E(n6406), .CP(clk), .QN(n27090) );
  EDFD1 \Mem_reg[74][13]  ( .D(n24749), .E(n6405), .CP(clk), .QN(n5709) );
  EDFD1 \Mem_reg[73][13]  ( .D(n24749), .E(n6404), .CP(clk), .QN(n27091) );
  EDFD1 \Mem_reg[72][13]  ( .D(n24749), .E(n6403), .CP(clk), .QN(n5613) );
  EDFD1 \Mem_reg[71][13]  ( .D(n24749), .E(n6402), .CP(clk), .QN(n5565) );
  EDFD1 \Mem_reg[70][13]  ( .D(n24749), .E(n6401), .CP(clk), .QN(n5517) );
  EDFD1 \Mem_reg[69][13]  ( .D(n24749), .E(n6400), .CP(clk), .QN(n5469) );
  EDFD1 \Mem_reg[68][13]  ( .D(n24749), .E(n6399), .CP(clk), .QN(n5421) );
  EDFD1 \Mem_reg[67][13]  ( .D(n24749), .E(n6398), .CP(clk), .QN(n5373) );
  EDFD1 \Mem_reg[66][13]  ( .D(n24749), .E(n6397), .CP(clk), .QN(n5325) );
  EDFD1 \Mem_reg[65][13]  ( .D(n24749), .E(n6396), .CP(clk), .QN(n15501) );
  EDFD1 \Mem_reg[64][13]  ( .D(n24749), .E(n6395), .CP(clk), .QN(n5229) );
  EDFD1 \Mem_reg[63][13]  ( .D(n24749), .E(n6456), .CP(clk), .QN(n5181) );
  EDFD1 \Mem_reg[62][13]  ( .D(n24749), .E(n6455), .CP(clk), .QN(n5133) );
  EDFD1 \Mem_reg[61][13]  ( .D(n24749), .E(n6454), .CP(clk), .QN(n17966) );
  EDFD1 \Mem_reg[60][13]  ( .D(n24749), .E(n6453), .CP(clk), .QN(n17965) );
  EDFD1 \Mem_reg[59][13]  ( .D(n24749), .E(n6452), .CP(clk), .QN(n4989) );
  EDFD1 \Mem_reg[58][13]  ( .D(n24749), .E(n6451), .CP(clk), .QN(n4941) );
  EDFD1 \Mem_reg[57][13]  ( .D(n24749), .E(n6450), .CP(clk), .QN(n4893) );
  EDFD1 \Mem_reg[56][13]  ( .D(n24749), .E(n6449), .CP(clk), .QN(n4845) );
  EDFD1 \Mem_reg[55][13]  ( .D(n24749), .E(n6448), .CP(clk), .QN(n4797) );
  EDFD1 \Mem_reg[54][13]  ( .D(n24749), .E(n6447), .CP(clk), .QN(n15500) );
  EDFD1 \Mem_reg[53][13]  ( .D(n24749), .E(n6446), .CP(clk), .QN(n4701) );
  EDFD1 \Mem_reg[52][13]  ( .D(n24749), .E(n6445), .CP(clk), .Q(n27088) );
  EDFD1 \Mem_reg[51][13]  ( .D(n24749), .E(n6444), .CP(clk), .QN(n4605) );
  EDFD1 \Mem_reg[50][13]  ( .D(n24749), .E(n6443), .CP(clk), .QN(n4557) );
  EDFD1 \Mem_reg[49][13]  ( .D(n24749), .E(n6442), .CP(clk), .QN(n4509) );
  EDFD1 \Mem_reg[48][13]  ( .D(n24749), .E(n6441), .CP(clk), .QN(n4461) );
  EDFD1 \Mem_reg[47][13]  ( .D(n24749), .E(n6440), .CP(clk), .QN(n4413) );
  EDFD1 \Mem_reg[46][13]  ( .D(n24749), .E(n6439), .CP(clk), .QN(n4365) );
  EDFD1 \Mem_reg[43][13]  ( .D(n24749), .E(n6438), .CP(clk), .QN(n4317) );
  EDFD1 \Mem_reg[42][13]  ( .D(n24749), .E(n6437), .CP(clk), .QN(n4269) );
  EDFD1 \Mem_reg[41][13]  ( .D(n24749), .E(n6436), .CP(clk), .QN(n4221) );
  EDFD1 \Mem_reg[40][13]  ( .D(n24749), .E(n6435), .CP(clk), .QN(n4173) );
  EDFD1 \Mem_reg[39][13]  ( .D(n24749), .E(n6434), .CP(clk), .QN(n4125) );
  EDFD1 \Mem_reg[38][13]  ( .D(n24749), .E(n6433), .CP(clk), .QN(n4077) );
  EDFD1 \Mem_reg[37][13]  ( .D(n24749), .E(n6432), .CP(clk), .QN(n4029) );
  EDFD1 \Mem_reg[36][13]  ( .D(n24749), .E(n6431), .CP(clk), .QN(n3981) );
  EDFD1 \Mem_reg[35][13]  ( .D(n24749), .E(n6430), .CP(clk), .QN(n3933) );
  EDFD1 \Mem_reg[34][13]  ( .D(n24749), .E(n6429), .CP(clk), .QN(n3885) );
  EDFD1 \Mem_reg[33][13]  ( .D(n24749), .E(n6428), .CP(clk), .QN(n3837) );
  EDFD1 \Mem_reg[32][13]  ( .D(n24749), .E(n6427), .CP(clk), .QN(n3789) );
  EDFD1 \Mem_reg[31][13]  ( .D(n24749), .E(n6426), .CP(clk), .QN(n3741) );
  EDFD1 \Mem_reg[30][13]  ( .D(n24749), .E(n6425), .CP(clk), .QN(n3693) );
  EDFD1 \Mem_reg[29][13]  ( .D(n24749), .E(n6424), .CP(clk), .QN(n3645) );
  EDFD1 \Mem_reg[28][13]  ( .D(n24749), .E(n6423), .CP(clk), .QN(n3597) );
  EDFD1 \Mem_reg[27][13]  ( .D(n24749), .E(n6422), .CP(clk), .QN(n3549) );
  EDFD1 \Mem_reg[26][13]  ( .D(n24749), .E(n6421), .CP(clk), .QN(n3501) );
  EDFD1 \Mem_reg[25][13]  ( .D(n24749), .E(n6420), .CP(clk), .QN(n3453) );
  EDFD1 \Mem_reg[24][13]  ( .D(n24749), .E(n6463), .CP(clk), .QN(n3405) );
  EDFD1 \Mem_reg[23][13]  ( .D(n24749), .E(n6464), .CP(clk), .QN(n3357) );
  EDFD1 \Mem_reg[22][13]  ( .D(n24749), .E(n6465), .CP(clk), .QN(n3309) );
  EDFD1 \Mem_reg[21][13]  ( .D(n24749), .E(n6466), .CP(clk), .QN(n3261) );
  EDFD1 \Mem_reg[20][13]  ( .D(n24749), .E(n6467), .CP(clk), .QN(n3213) );
  EDFD1 \Mem_reg[19][13]  ( .D(n24749), .E(n6468), .CP(clk), .QN(n3165) );
  EDFD1 \Mem_reg[18][13]  ( .D(n24749), .E(n6469), .CP(clk), .QN(n3117) );
  EDFD1 \Mem_reg[17][13]  ( .D(n24749), .E(n6470), .CP(clk), .QN(n3069) );
  EDFD1 \Mem_reg[16][13]  ( .D(n24749), .E(n6471), .CP(clk), .QN(n3021) );
  EDFD1 \Mem_reg[15][13]  ( .D(n24749), .E(n6472), .CP(clk), .QN(n2973) );
  EDFD1 \Mem_reg[14][13]  ( .D(n24749), .E(n24720), .CP(clk), .QN(n2925) );
  EDFD1 \Mem_reg[13][13]  ( .D(n24749), .E(n24709), .CP(clk), .QN(n2877) );
  EDFD1 \Mem_reg[12][13]  ( .D(n24749), .E(n24717), .CP(clk), .QN(n2829) );
  EDFD1 \Mem_reg[11][13]  ( .D(n24749), .E(n24707), .CP(clk), .QN(n2781) );
  EDFD1 \Mem_reg[10][13]  ( .D(n24749), .E(n6477), .CP(clk), .QN(n2733) );
  EDFD1 \Mem_reg[9][13]  ( .D(n24749), .E(n24708), .CP(clk), .QN(n2685) );
  EDFD1 \Mem_reg[8][13]  ( .D(n24749), .E(n15642), .CP(clk), .QN(n2637) );
  EDFD1 \Mem_reg[7][13]  ( .D(n24749), .E(n24718), .CP(clk), .QN(n2589) );
  EDFD1 \Mem_reg[6][13]  ( .D(n24749), .E(n24716), .CP(clk), .QN(n2541) );
  EDFD1 \Mem_reg[5][13]  ( .D(n24749), .E(n24719), .CP(clk), .QN(n2493) );
  EDFD1 \Mem_reg[4][13]  ( .D(n24749), .E(n24706), .CP(clk), .QN(n2445) );
  EDFD1 \Mem_reg[3][13]  ( .D(n24749), .E(n24721), .CP(clk), .QN(n2397) );
  EDFD1 \Mem_reg[2][13]  ( .D(n24749), .E(n6460), .CP(clk), .QN(n2349) );
  EDFD1 \Mem_reg[1][13]  ( .D(n24749), .E(n24703), .CP(clk), .QN(n2301) );
  EDFD1 \Mem_reg[0][13]  ( .D(n24749), .E(n24705), .CP(clk), .QN(n2253) );
  EDFD1 \Mem_reg[88][12]  ( .D(n24747), .E(n6419), .CP(clk), .Q(n27085) );
  EDFD1 \Mem_reg[87][12]  ( .D(n24747), .E(n6418), .CP(clk), .QN(n6334) );
  EDFD1 \Mem_reg[86][12]  ( .D(n24747), .E(n6417), .CP(clk), .QN(n24595) );
  EDFD1 \Mem_reg[85][12]  ( .D(n24747), .E(n6416), .CP(clk), .QN(n6238) );
  EDFD1 \Mem_reg[84][12]  ( .D(n24747), .E(n6415), .CP(clk), .QN(n6190) );
  EDFD1 \Mem_reg[83][12]  ( .D(n24747), .E(n6414), .CP(clk), .QN(n6142) );
  EDFD1 \Mem_reg[82][12]  ( .D(n24747), .E(n6413), .CP(clk), .QN(n6094) );
  EDFD1 \Mem_reg[81][12]  ( .D(n24747), .E(n6412), .CP(clk), .QN(n6046) );
  EDFD1 \Mem_reg[80][12]  ( .D(n24747), .E(n6411), .CP(clk), .QN(n5998) );
  EDFD1 \Mem_reg[79][12]  ( .D(n24747), .E(n6410), .CP(clk), .QN(n5950) );
  EDFD1 \Mem_reg[78][12]  ( .D(n24747), .E(n6409), .CP(clk), .QN(n5902) );
  EDFD1 \Mem_reg[77][12]  ( .D(n24747), .E(n6408), .CP(clk), .QN(n5854) );
  EDFD1 \Mem_reg[76][12]  ( .D(n24747), .E(n6407), .CP(clk), .QN(n5806) );
  EDFD1 \Mem_reg[75][12]  ( .D(n24747), .E(n6406), .CP(clk), .QN(n27086) );
  EDFD1 \Mem_reg[74][12]  ( .D(n24747), .E(n6405), .CP(clk), .QN(n5710) );
  EDFD1 \Mem_reg[73][12]  ( .D(n24747), .E(n6404), .CP(clk), .QN(n27087) );
  EDFD1 \Mem_reg[72][12]  ( .D(n24747), .E(n6403), .CP(clk), .QN(n5614) );
  EDFD1 \Mem_reg[71][12]  ( .D(n24747), .E(n6402), .CP(clk), .QN(n5566) );
  EDFD1 \Mem_reg[70][12]  ( .D(n24747), .E(n6401), .CP(clk), .QN(n5518) );
  EDFD1 \Mem_reg[69][12]  ( .D(n24747), .E(n6400), .CP(clk), .QN(n5470) );
  EDFD1 \Mem_reg[68][12]  ( .D(n24747), .E(n6399), .CP(clk), .QN(n5422) );
  EDFD1 \Mem_reg[67][12]  ( .D(n24747), .E(n6398), .CP(clk), .QN(n5374) );
  EDFD1 \Mem_reg[66][12]  ( .D(n24747), .E(n6397), .CP(clk), .QN(n5326) );
  EDFD1 \Mem_reg[65][12]  ( .D(n24747), .E(n6396), .CP(clk), .QN(n15497) );
  EDFD1 \Mem_reg[64][12]  ( .D(n24747), .E(n6395), .CP(clk), .QN(n5230) );
  EDFD1 \Mem_reg[63][12]  ( .D(n24747), .E(n6456), .CP(clk), .QN(n5182) );
  EDFD1 \Mem_reg[62][12]  ( .D(n24747), .E(n6455), .CP(clk), .QN(n5134) );
  EDFD1 \Mem_reg[61][12]  ( .D(n24747), .E(n6454), .CP(clk), .QN(n17963) );
  EDFD1 \Mem_reg[60][12]  ( .D(n24747), .E(n6453), .CP(clk), .QN(n17962) );
  EDFD1 \Mem_reg[59][12]  ( .D(n24747), .E(n6452), .CP(clk), .QN(n4990) );
  EDFD1 \Mem_reg[58][12]  ( .D(n24747), .E(n6451), .CP(clk), .QN(n4942) );
  EDFD1 \Mem_reg[57][12]  ( .D(n24747), .E(n6450), .CP(clk), .QN(n4894) );
  EDFD1 \Mem_reg[56][12]  ( .D(n24747), .E(n6449), .CP(clk), .QN(n4846) );
  EDFD1 \Mem_reg[55][12]  ( .D(n24747), .E(n6448), .CP(clk), .QN(n4798) );
  EDFD1 \Mem_reg[54][12]  ( .D(n24747), .E(n6447), .CP(clk), .QN(n15496) );
  EDFD1 \Mem_reg[53][12]  ( .D(n24747), .E(n6446), .CP(clk), .QN(n4702) );
  EDFD1 \Mem_reg[52][12]  ( .D(n24747), .E(n6445), .CP(clk), .Q(n27084) );
  EDFD1 \Mem_reg[51][12]  ( .D(n24747), .E(n6444), .CP(clk), .QN(n4606) );
  EDFD1 \Mem_reg[50][12]  ( .D(n24747), .E(n6443), .CP(clk), .QN(n4558) );
  EDFD1 \Mem_reg[49][12]  ( .D(n24747), .E(n6442), .CP(clk), .QN(n4510) );
  EDFD1 \Mem_reg[48][12]  ( .D(n24747), .E(n6441), .CP(clk), .QN(n4462) );
  EDFD1 \Mem_reg[47][12]  ( .D(n24747), .E(n6440), .CP(clk), .QN(n4414) );
  EDFD1 \Mem_reg[46][12]  ( .D(n24747), .E(n6439), .CP(clk), .QN(n4366) );
  EDFD1 \Mem_reg[43][12]  ( .D(n24747), .E(n6438), .CP(clk), .QN(n4318) );
  EDFD1 \Mem_reg[42][12]  ( .D(n24747), .E(n6437), .CP(clk), .QN(n4270) );
  EDFD1 \Mem_reg[41][12]  ( .D(n24747), .E(n6436), .CP(clk), .QN(n4222) );
  EDFD1 \Mem_reg[40][12]  ( .D(n24747), .E(n6435), .CP(clk), .QN(n4174) );
  EDFD1 \Mem_reg[39][12]  ( .D(n24747), .E(n6434), .CP(clk), .QN(n4126) );
  EDFD1 \Mem_reg[38][12]  ( .D(n24747), .E(n6433), .CP(clk), .QN(n4078) );
  EDFD1 \Mem_reg[37][12]  ( .D(n24747), .E(n6432), .CP(clk), .QN(n4030) );
  EDFD1 \Mem_reg[36][12]  ( .D(n24747), .E(n6431), .CP(clk), .QN(n3982) );
  EDFD1 \Mem_reg[35][12]  ( .D(n24747), .E(n6430), .CP(clk), .QN(n3934) );
  EDFD1 \Mem_reg[34][12]  ( .D(n24747), .E(n6429), .CP(clk), .QN(n3886) );
  EDFD1 \Mem_reg[33][12]  ( .D(n24747), .E(n6428), .CP(clk), .QN(n3838) );
  EDFD1 \Mem_reg[32][12]  ( .D(n24747), .E(n6427), .CP(clk), .QN(n3790) );
  EDFD1 \Mem_reg[31][12]  ( .D(n24747), .E(n6426), .CP(clk), .QN(n3742) );
  EDFD1 \Mem_reg[30][12]  ( .D(n24747), .E(n6425), .CP(clk), .QN(n3694) );
  EDFD1 \Mem_reg[29][12]  ( .D(n24747), .E(n6424), .CP(clk), .QN(n3646) );
  EDFD1 \Mem_reg[28][12]  ( .D(n24747), .E(n6423), .CP(clk), .QN(n3598) );
  EDFD1 \Mem_reg[27][12]  ( .D(n24747), .E(n6422), .CP(clk), .QN(n3550) );
  EDFD1 \Mem_reg[26][12]  ( .D(n24747), .E(n6421), .CP(clk), .QN(n3502) );
  EDFD1 \Mem_reg[25][12]  ( .D(n24747), .E(n6420), .CP(clk), .QN(n3454) );
  EDFD1 \Mem_reg[24][12]  ( .D(n24747), .E(n6463), .CP(clk), .QN(n3406) );
  EDFD1 \Mem_reg[23][12]  ( .D(n24747), .E(n6464), .CP(clk), .QN(n3358) );
  EDFD1 \Mem_reg[22][12]  ( .D(n24747), .E(n6465), .CP(clk), .QN(n3310) );
  EDFD1 \Mem_reg[21][12]  ( .D(n24747), .E(n6466), .CP(clk), .QN(n3262) );
  EDFD1 \Mem_reg[20][12]  ( .D(n24747), .E(n6467), .CP(clk), .QN(n3214) );
  EDFD1 \Mem_reg[19][12]  ( .D(n24747), .E(n6468), .CP(clk), .QN(n3166) );
  EDFD1 \Mem_reg[18][12]  ( .D(n24747), .E(n6469), .CP(clk), .QN(n3118) );
  EDFD1 \Mem_reg[17][12]  ( .D(n24747), .E(n6470), .CP(clk), .QN(n3070) );
  EDFD1 \Mem_reg[16][12]  ( .D(n24747), .E(n6471), .CP(clk), .QN(n3022) );
  EDFD1 \Mem_reg[15][12]  ( .D(n24747), .E(n6472), .CP(clk), .QN(n2974) );
  EDFD1 \Mem_reg[14][12]  ( .D(n24747), .E(n24720), .CP(clk), .QN(n2926) );
  EDFD1 \Mem_reg[13][12]  ( .D(n24747), .E(n24709), .CP(clk), .QN(n2878) );
  EDFD1 \Mem_reg[12][12]  ( .D(n24747), .E(n24717), .CP(clk), .QN(n2830) );
  EDFD1 \Mem_reg[11][12]  ( .D(n24747), .E(n24707), .CP(clk), .QN(n2782) );
  EDFD1 \Mem_reg[10][12]  ( .D(n24747), .E(n6477), .CP(clk), .QN(n2734) );
  EDFD1 \Mem_reg[9][12]  ( .D(n24747), .E(n24708), .CP(clk), .QN(n2686) );
  EDFD1 \Mem_reg[8][12]  ( .D(n24747), .E(n15642), .CP(clk), .QN(n2638) );
  EDFD1 \Mem_reg[7][12]  ( .D(n24747), .E(n24718), .CP(clk), .QN(n2590) );
  EDFD1 \Mem_reg[6][12]  ( .D(n24747), .E(n24716), .CP(clk), .QN(n2542) );
  EDFD1 \Mem_reg[5][12]  ( .D(n24747), .E(n24719), .CP(clk), .QN(n2494) );
  EDFD1 \Mem_reg[4][12]  ( .D(n24747), .E(n24706), .CP(clk), .QN(n2446) );
  EDFD1 \Mem_reg[3][12]  ( .D(n24747), .E(n24721), .CP(clk), .QN(n2398) );
  EDFD1 \Mem_reg[2][12]  ( .D(n24747), .E(n6460), .CP(clk), .QN(n2350) );
  EDFD1 \Mem_reg[1][12]  ( .D(n24747), .E(n24703), .CP(clk), .QN(n2302) );
  EDFD1 \Mem_reg[0][12]  ( .D(n24747), .E(n24705), .CP(clk), .QN(n2254) );
  EDFD1 \Mem_reg[88][11]  ( .D(n24745), .E(n6419), .CP(clk), .Q(n27081) );
  EDFD1 \Mem_reg[87][11]  ( .D(n24745), .E(n6418), .CP(clk), .QN(n6335) );
  EDFD1 \Mem_reg[86][11]  ( .D(n24745), .E(n6417), .CP(clk), .QN(n24592) );
  EDFD1 \Mem_reg[85][11]  ( .D(n24745), .E(n6416), .CP(clk), .QN(n6239) );
  EDFD1 \Mem_reg[84][11]  ( .D(n24745), .E(n6415), .CP(clk), .QN(n6191) );
  EDFD1 \Mem_reg[83][11]  ( .D(n24745), .E(n6414), .CP(clk), .QN(n6143) );
  EDFD1 \Mem_reg[82][11]  ( .D(n24745), .E(n6413), .CP(clk), .QN(n6095) );
  EDFD1 \Mem_reg[81][11]  ( .D(n24745), .E(n6412), .CP(clk), .QN(n6047) );
  EDFD1 \Mem_reg[80][11]  ( .D(n24745), .E(n6411), .CP(clk), .QN(n5999) );
  EDFD1 \Mem_reg[79][11]  ( .D(n24745), .E(n6410), .CP(clk), .QN(n5951) );
  EDFD1 \Mem_reg[78][11]  ( .D(n24745), .E(n6409), .CP(clk), .QN(n5903) );
  EDFD1 \Mem_reg[77][11]  ( .D(n24745), .E(n6408), .CP(clk), .QN(n5855) );
  EDFD1 \Mem_reg[76][11]  ( .D(n24745), .E(n6407), .CP(clk), .QN(n5807) );
  EDFD1 \Mem_reg[75][11]  ( .D(n24745), .E(n6406), .CP(clk), .QN(n27082) );
  EDFD1 \Mem_reg[74][11]  ( .D(n24745), .E(n6405), .CP(clk), .QN(n5711) );
  EDFD1 \Mem_reg[73][11]  ( .D(n24745), .E(n6404), .CP(clk), .QN(n27083) );
  EDFD1 \Mem_reg[72][11]  ( .D(n24745), .E(n6403), .CP(clk), .QN(n5615) );
  EDFD1 \Mem_reg[71][11]  ( .D(n24745), .E(n6402), .CP(clk), .QN(n5567) );
  EDFD1 \Mem_reg[70][11]  ( .D(n24745), .E(n6401), .CP(clk), .QN(n5519) );
  EDFD1 \Mem_reg[69][11]  ( .D(n24745), .E(n6400), .CP(clk), .QN(n5471) );
  EDFD1 \Mem_reg[68][11]  ( .D(n24745), .E(n6399), .CP(clk), .QN(n5423) );
  EDFD1 \Mem_reg[67][11]  ( .D(n24745), .E(n6398), .CP(clk), .QN(n5375) );
  EDFD1 \Mem_reg[66][11]  ( .D(n24745), .E(n6397), .CP(clk), .QN(n5327) );
  EDFD1 \Mem_reg[65][11]  ( .D(n24745), .E(n6396), .CP(clk), .QN(n15493) );
  EDFD1 \Mem_reg[64][11]  ( .D(n24745), .E(n6395), .CP(clk), .QN(n5231) );
  EDFD1 \Mem_reg[63][11]  ( .D(n24745), .E(n6456), .CP(clk), .QN(n5183) );
  EDFD1 \Mem_reg[62][11]  ( .D(n24745), .E(n6455), .CP(clk), .QN(n5135) );
  EDFD1 \Mem_reg[61][11]  ( .D(n24745), .E(n6454), .CP(clk), .QN(n17960) );
  EDFD1 \Mem_reg[60][11]  ( .D(n24745), .E(n6453), .CP(clk), .QN(n17959) );
  EDFD1 \Mem_reg[59][11]  ( .D(n24745), .E(n6452), .CP(clk), .QN(n4991) );
  EDFD1 \Mem_reg[58][11]  ( .D(n24745), .E(n6451), .CP(clk), .QN(n4943) );
  EDFD1 \Mem_reg[57][11]  ( .D(n24745), .E(n6450), .CP(clk), .QN(n4895) );
  EDFD1 \Mem_reg[56][11]  ( .D(n24745), .E(n6449), .CP(clk), .QN(n4847) );
  EDFD1 \Mem_reg[55][11]  ( .D(n24745), .E(n6448), .CP(clk), .QN(n4799) );
  EDFD1 \Mem_reg[54][11]  ( .D(n24745), .E(n6447), .CP(clk), .QN(n15492) );
  EDFD1 \Mem_reg[53][11]  ( .D(n24745), .E(n6446), .CP(clk), .QN(n4703) );
  EDFD1 \Mem_reg[52][11]  ( .D(n24745), .E(n6445), .CP(clk), .Q(n27080) );
  EDFD1 \Mem_reg[51][11]  ( .D(n24745), .E(n6444), .CP(clk), .QN(n4607) );
  EDFD1 \Mem_reg[50][11]  ( .D(n24745), .E(n6443), .CP(clk), .QN(n4559) );
  EDFD1 \Mem_reg[49][11]  ( .D(n24745), .E(n6442), .CP(clk), .QN(n4511) );
  EDFD1 \Mem_reg[48][11]  ( .D(n24745), .E(n6441), .CP(clk), .QN(n4463) );
  EDFD1 \Mem_reg[47][11]  ( .D(n24745), .E(n6440), .CP(clk), .QN(n4415) );
  EDFD1 \Mem_reg[46][11]  ( .D(n24745), .E(n6439), .CP(clk), .QN(n4367) );
  EDFD1 \Mem_reg[43][11]  ( .D(n24745), .E(n6438), .CP(clk), .QN(n4319) );
  EDFD1 \Mem_reg[42][11]  ( .D(n24745), .E(n6437), .CP(clk), .QN(n4271) );
  EDFD1 \Mem_reg[41][11]  ( .D(n24745), .E(n6436), .CP(clk), .QN(n4223) );
  EDFD1 \Mem_reg[40][11]  ( .D(n24745), .E(n6435), .CP(clk), .QN(n4175) );
  EDFD1 \Mem_reg[39][11]  ( .D(n24745), .E(n6434), .CP(clk), .QN(n4127) );
  EDFD1 \Mem_reg[38][11]  ( .D(n24745), .E(n6433), .CP(clk), .QN(n4079) );
  EDFD1 \Mem_reg[37][11]  ( .D(n24745), .E(n6432), .CP(clk), .QN(n4031) );
  EDFD1 \Mem_reg[36][11]  ( .D(n24745), .E(n6431), .CP(clk), .QN(n3983) );
  EDFD1 \Mem_reg[35][11]  ( .D(n24745), .E(n6430), .CP(clk), .QN(n3935) );
  EDFD1 \Mem_reg[34][11]  ( .D(n24745), .E(n6429), .CP(clk), .QN(n3887) );
  EDFD1 \Mem_reg[33][11]  ( .D(n24745), .E(n6428), .CP(clk), .QN(n3839) );
  EDFD1 \Mem_reg[32][11]  ( .D(n24745), .E(n6427), .CP(clk), .QN(n3791) );
  EDFD1 \Mem_reg[31][11]  ( .D(n24745), .E(n6426), .CP(clk), .QN(n3743) );
  EDFD1 \Mem_reg[30][11]  ( .D(n24745), .E(n6425), .CP(clk), .QN(n3695) );
  EDFD1 \Mem_reg[29][11]  ( .D(n24745), .E(n6424), .CP(clk), .QN(n3647) );
  EDFD1 \Mem_reg[28][11]  ( .D(n24745), .E(n6423), .CP(clk), .QN(n3599) );
  EDFD1 \Mem_reg[27][11]  ( .D(n24745), .E(n6422), .CP(clk), .QN(n3551) );
  EDFD1 \Mem_reg[26][11]  ( .D(n24745), .E(n6421), .CP(clk), .QN(n3503) );
  EDFD1 \Mem_reg[25][11]  ( .D(n24745), .E(n6420), .CP(clk), .QN(n3455) );
  EDFD1 \Mem_reg[24][11]  ( .D(n24745), .E(n6463), .CP(clk), .QN(n3407) );
  EDFD1 \Mem_reg[23][11]  ( .D(n24745), .E(n6464), .CP(clk), .QN(n3359) );
  EDFD1 \Mem_reg[22][11]  ( .D(n24745), .E(n6465), .CP(clk), .QN(n3311) );
  EDFD1 \Mem_reg[21][11]  ( .D(n24745), .E(n6466), .CP(clk), .QN(n3263) );
  EDFD1 \Mem_reg[20][11]  ( .D(n24745), .E(n6467), .CP(clk), .QN(n3215) );
  EDFD1 \Mem_reg[19][11]  ( .D(n24745), .E(n6468), .CP(clk), .QN(n3167) );
  EDFD1 \Mem_reg[18][11]  ( .D(n24745), .E(n6469), .CP(clk), .QN(n3119) );
  EDFD1 \Mem_reg[17][11]  ( .D(n24745), .E(n6470), .CP(clk), .QN(n3071) );
  EDFD1 \Mem_reg[16][11]  ( .D(n24745), .E(n6471), .CP(clk), .QN(n3023) );
  EDFD1 \Mem_reg[15][11]  ( .D(n24745), .E(n6472), .CP(clk), .QN(n2975) );
  EDFD1 \Mem_reg[14][11]  ( .D(n24745), .E(n24720), .CP(clk), .QN(n2927) );
  EDFD1 \Mem_reg[13][11]  ( .D(n24745), .E(n24709), .CP(clk), .QN(n2879) );
  EDFD1 \Mem_reg[12][11]  ( .D(n24745), .E(n24717), .CP(clk), .QN(n2831) );
  EDFD1 \Mem_reg[11][11]  ( .D(n24745), .E(n24707), .CP(clk), .QN(n2783) );
  EDFD1 \Mem_reg[10][11]  ( .D(n24745), .E(n6477), .CP(clk), .QN(n2735) );
  EDFD1 \Mem_reg[9][11]  ( .D(n24745), .E(n24708), .CP(clk), .QN(n2687) );
  EDFD1 \Mem_reg[8][11]  ( .D(n24745), .E(n15642), .CP(clk), .QN(n2639) );
  EDFD1 \Mem_reg[7][11]  ( .D(n24745), .E(n24718), .CP(clk), .QN(n2591) );
  EDFD1 \Mem_reg[6][11]  ( .D(n24745), .E(n24716), .CP(clk), .QN(n2543) );
  EDFD1 \Mem_reg[5][11]  ( .D(n24745), .E(n24719), .CP(clk), .QN(n2495) );
  EDFD1 \Mem_reg[4][11]  ( .D(n24745), .E(n24706), .CP(clk), .QN(n2447) );
  EDFD1 \Mem_reg[3][11]  ( .D(n24745), .E(n24721), .CP(clk), .QN(n2399) );
  EDFD1 \Mem_reg[2][11]  ( .D(n24745), .E(n6460), .CP(clk), .QN(n2351) );
  EDFD1 \Mem_reg[1][11]  ( .D(n24745), .E(n24703), .CP(clk), .QN(n2303) );
  EDFD1 \Mem_reg[0][11]  ( .D(n24745), .E(n24705), .CP(clk), .QN(n2255) );
  EDFD1 \Mem_reg[88][10]  ( .D(n24743), .E(n6419), .CP(clk), .Q(n27077) );
  EDFD1 \Mem_reg[87][10]  ( .D(n24743), .E(n6418), .CP(clk), .QN(n6336) );
  EDFD1 \Mem_reg[86][10]  ( .D(n24743), .E(n6417), .CP(clk), .QN(n24589) );
  EDFD1 \Mem_reg[85][10]  ( .D(n24743), .E(n6416), .CP(clk), .QN(n6240) );
  EDFD1 \Mem_reg[84][10]  ( .D(n24743), .E(n6415), .CP(clk), .QN(n6192) );
  EDFD1 \Mem_reg[83][10]  ( .D(n24743), .E(n6414), .CP(clk), .QN(n6144) );
  EDFD1 \Mem_reg[82][10]  ( .D(n24743), .E(n6413), .CP(clk), .QN(n6096) );
  EDFD1 \Mem_reg[81][10]  ( .D(n24743), .E(n6412), .CP(clk), .QN(n6048) );
  EDFD1 \Mem_reg[80][10]  ( .D(n24743), .E(n6411), .CP(clk), .QN(n6000) );
  EDFD1 \Mem_reg[79][10]  ( .D(n24743), .E(n6410), .CP(clk), .QN(n5952) );
  EDFD1 \Mem_reg[78][10]  ( .D(n24743), .E(n6409), .CP(clk), .QN(n5904) );
  EDFD1 \Mem_reg[77][10]  ( .D(n24743), .E(n6408), .CP(clk), .QN(n5856) );
  EDFD1 \Mem_reg[76][10]  ( .D(n24743), .E(n6407), .CP(clk), .QN(n5808) );
  EDFD1 \Mem_reg[75][10]  ( .D(n24743), .E(n6406), .CP(clk), .QN(n27078) );
  EDFD1 \Mem_reg[74][10]  ( .D(n24743), .E(n6405), .CP(clk), .QN(n5712) );
  EDFD1 \Mem_reg[73][10]  ( .D(n24743), .E(n6404), .CP(clk), .QN(n27079) );
  EDFD1 \Mem_reg[72][10]  ( .D(n24743), .E(n6403), .CP(clk), .QN(n5616) );
  EDFD1 \Mem_reg[71][10]  ( .D(n24743), .E(n6402), .CP(clk), .QN(n5568) );
  EDFD1 \Mem_reg[70][10]  ( .D(n24743), .E(n6401), .CP(clk), .QN(n5520) );
  EDFD1 \Mem_reg[69][10]  ( .D(n24743), .E(n6400), .CP(clk), .QN(n5472) );
  EDFD1 \Mem_reg[68][10]  ( .D(n24743), .E(n6399), .CP(clk), .QN(n5424) );
  EDFD1 \Mem_reg[67][10]  ( .D(n24743), .E(n6398), .CP(clk), .QN(n5376) );
  EDFD1 \Mem_reg[66][10]  ( .D(n24743), .E(n6397), .CP(clk), .QN(n5328) );
  EDFD1 \Mem_reg[65][10]  ( .D(n24743), .E(n6396), .CP(clk), .QN(n15489) );
  EDFD1 \Mem_reg[64][10]  ( .D(n24743), .E(n6395), .CP(clk), .QN(n5232) );
  EDFD1 \Mem_reg[63][10]  ( .D(n24743), .E(n6456), .CP(clk), .QN(n5184) );
  EDFD1 \Mem_reg[62][10]  ( .D(n24743), .E(n6455), .CP(clk), .QN(n5136) );
  EDFD1 \Mem_reg[61][10]  ( .D(n24743), .E(n6454), .CP(clk), .QN(n17957) );
  EDFD1 \Mem_reg[60][10]  ( .D(n24743), .E(n6453), .CP(clk), .QN(n17956) );
  EDFD1 \Mem_reg[59][10]  ( .D(n24743), .E(n6452), .CP(clk), .QN(n4992) );
  EDFD1 \Mem_reg[58][10]  ( .D(n24743), .E(n6451), .CP(clk), .QN(n4944) );
  EDFD1 \Mem_reg[57][10]  ( .D(n24743), .E(n6450), .CP(clk), .QN(n4896) );
  EDFD1 \Mem_reg[56][10]  ( .D(n24743), .E(n6449), .CP(clk), .QN(n4848) );
  EDFD1 \Mem_reg[55][10]  ( .D(n24743), .E(n6448), .CP(clk), .QN(n4800) );
  EDFD1 \Mem_reg[54][10]  ( .D(n24743), .E(n6447), .CP(clk), .QN(n15488) );
  EDFD1 \Mem_reg[53][10]  ( .D(n24743), .E(n6446), .CP(clk), .QN(n4704) );
  EDFD1 \Mem_reg[52][10]  ( .D(n24743), .E(n6445), .CP(clk), .Q(n27076) );
  EDFD1 \Mem_reg[51][10]  ( .D(n24743), .E(n6444), .CP(clk), .QN(n4608) );
  EDFD1 \Mem_reg[50][10]  ( .D(n24743), .E(n6443), .CP(clk), .QN(n4560) );
  EDFD1 \Mem_reg[49][10]  ( .D(n24743), .E(n6442), .CP(clk), .QN(n4512) );
  EDFD1 \Mem_reg[48][10]  ( .D(n24743), .E(n6441), .CP(clk), .QN(n4464) );
  EDFD1 \Mem_reg[47][10]  ( .D(n24743), .E(n6440), .CP(clk), .QN(n4416) );
  EDFD1 \Mem_reg[46][10]  ( .D(n24743), .E(n6439), .CP(clk), .QN(n4368) );
  EDFD1 \Mem_reg[43][10]  ( .D(n24743), .E(n6438), .CP(clk), .QN(n4320) );
  EDFD1 \Mem_reg[42][10]  ( .D(n24743), .E(n6437), .CP(clk), .QN(n4272) );
  EDFD1 \Mem_reg[41][10]  ( .D(n24743), .E(n6436), .CP(clk), .QN(n4224) );
  EDFD1 \Mem_reg[40][10]  ( .D(n24743), .E(n6435), .CP(clk), .QN(n4176) );
  EDFD1 \Mem_reg[39][10]  ( .D(n24743), .E(n6434), .CP(clk), .QN(n4128) );
  EDFD1 \Mem_reg[38][10]  ( .D(n24743), .E(n6433), .CP(clk), .QN(n4080) );
  EDFD1 \Mem_reg[37][10]  ( .D(n24743), .E(n6432), .CP(clk), .QN(n4032) );
  EDFD1 \Mem_reg[36][10]  ( .D(n24743), .E(n6431), .CP(clk), .QN(n3984) );
  EDFD1 \Mem_reg[35][10]  ( .D(n24743), .E(n6430), .CP(clk), .QN(n3936) );
  EDFD1 \Mem_reg[34][10]  ( .D(n24743), .E(n6429), .CP(clk), .QN(n3888) );
  EDFD1 \Mem_reg[33][10]  ( .D(n24743), .E(n6428), .CP(clk), .QN(n3840) );
  EDFD1 \Mem_reg[32][10]  ( .D(n24743), .E(n6427), .CP(clk), .QN(n3792) );
  EDFD1 \Mem_reg[31][10]  ( .D(n24743), .E(n6426), .CP(clk), .QN(n3744) );
  EDFD1 \Mem_reg[30][10]  ( .D(n24743), .E(n6425), .CP(clk), .QN(n3696) );
  EDFD1 \Mem_reg[29][10]  ( .D(n24743), .E(n6424), .CP(clk), .QN(n3648) );
  EDFD1 \Mem_reg[28][10]  ( .D(n24743), .E(n6423), .CP(clk), .QN(n3600) );
  EDFD1 \Mem_reg[27][10]  ( .D(n24743), .E(n6422), .CP(clk), .QN(n3552) );
  EDFD1 \Mem_reg[26][10]  ( .D(n24743), .E(n6421), .CP(clk), .QN(n3504) );
  EDFD1 \Mem_reg[25][10]  ( .D(n24743), .E(n6420), .CP(clk), .QN(n3456) );
  EDFD1 \Mem_reg[24][10]  ( .D(n24743), .E(n6463), .CP(clk), .QN(n3408) );
  EDFD1 \Mem_reg[23][10]  ( .D(n24743), .E(n6464), .CP(clk), .QN(n3360) );
  EDFD1 \Mem_reg[22][10]  ( .D(n24743), .E(n6465), .CP(clk), .QN(n3312) );
  EDFD1 \Mem_reg[21][10]  ( .D(n24743), .E(n6466), .CP(clk), .QN(n3264) );
  EDFD1 \Mem_reg[20][10]  ( .D(n24743), .E(n6467), .CP(clk), .QN(n3216) );
  EDFD1 \Mem_reg[19][10]  ( .D(n24743), .E(n6468), .CP(clk), .QN(n3168) );
  EDFD1 \Mem_reg[18][10]  ( .D(n24743), .E(n6469), .CP(clk), .QN(n3120) );
  EDFD1 \Mem_reg[17][10]  ( .D(n24743), .E(n6470), .CP(clk), .QN(n3072) );
  EDFD1 \Mem_reg[16][10]  ( .D(n24743), .E(n6471), .CP(clk), .QN(n3024) );
  EDFD1 \Mem_reg[15][10]  ( .D(n24743), .E(n6472), .CP(clk), .QN(n2976) );
  EDFD1 \Mem_reg[14][10]  ( .D(n24743), .E(n24720), .CP(clk), .QN(n2928) );
  EDFD1 \Mem_reg[13][10]  ( .D(n24743), .E(n24709), .CP(clk), .QN(n2880) );
  EDFD1 \Mem_reg[12][10]  ( .D(n24743), .E(n24717), .CP(clk), .QN(n2832) );
  EDFD1 \Mem_reg[11][10]  ( .D(n24743), .E(n24707), .CP(clk), .QN(n2784) );
  EDFD1 \Mem_reg[10][10]  ( .D(n24743), .E(n6477), .CP(clk), .QN(n2736) );
  EDFD1 \Mem_reg[9][10]  ( .D(n24743), .E(n24708), .CP(clk), .QN(n2688) );
  EDFD1 \Mem_reg[8][10]  ( .D(n24743), .E(n15642), .CP(clk), .QN(n2640) );
  EDFD1 \Mem_reg[7][10]  ( .D(n24743), .E(n24718), .CP(clk), .QN(n2592) );
  EDFD1 \Mem_reg[6][10]  ( .D(n24743), .E(n24716), .CP(clk), .QN(n2544) );
  EDFD1 \Mem_reg[5][10]  ( .D(n24743), .E(n24719), .CP(clk), .QN(n2496) );
  EDFD1 \Mem_reg[4][10]  ( .D(n24743), .E(n24706), .CP(clk), .QN(n2448) );
  EDFD1 \Mem_reg[3][10]  ( .D(n24743), .E(n24721), .CP(clk), .QN(n2400) );
  EDFD1 \Mem_reg[2][10]  ( .D(n24743), .E(n6460), .CP(clk), .QN(n2352) );
  EDFD1 \Mem_reg[1][10]  ( .D(n24743), .E(n24703), .CP(clk), .QN(n2304) );
  EDFD1 \Mem_reg[0][10]  ( .D(n24743), .E(n24705), .CP(clk), .QN(n2256) );
  EDFD1 \Mem_reg[88][9]  ( .D(n24741), .E(n6419), .CP(clk), .Q(n27073) );
  EDFD1 \Mem_reg[87][9]  ( .D(n24741), .E(n6418), .CP(clk), .QN(n6337) );
  EDFD1 \Mem_reg[86][9]  ( .D(n24741), .E(n6417), .CP(clk), .QN(n24586) );
  EDFD1 \Mem_reg[85][9]  ( .D(n24741), .E(n6416), .CP(clk), .QN(n6241) );
  EDFD1 \Mem_reg[84][9]  ( .D(n24741), .E(n6415), .CP(clk), .QN(n6193) );
  EDFD1 \Mem_reg[83][9]  ( .D(n24741), .E(n6414), .CP(clk), .QN(n6145) );
  EDFD1 \Mem_reg[82][9]  ( .D(n24741), .E(n6413), .CP(clk), .QN(n6097) );
  EDFD1 \Mem_reg[81][9]  ( .D(n24741), .E(n6412), .CP(clk), .QN(n6049) );
  EDFD1 \Mem_reg[80][9]  ( .D(n24741), .E(n6411), .CP(clk), .QN(n6001) );
  EDFD1 \Mem_reg[79][9]  ( .D(n24741), .E(n6410), .CP(clk), .QN(n5953) );
  EDFD1 \Mem_reg[78][9]  ( .D(n24741), .E(n6409), .CP(clk), .QN(n5905) );
  EDFD1 \Mem_reg[77][9]  ( .D(n24741), .E(n6408), .CP(clk), .QN(n5857) );
  EDFD1 \Mem_reg[76][9]  ( .D(n24741), .E(n6407), .CP(clk), .QN(n5809) );
  EDFD1 \Mem_reg[75][9]  ( .D(n24741), .E(n6406), .CP(clk), .QN(n27074) );
  EDFD1 \Mem_reg[74][9]  ( .D(n24741), .E(n6405), .CP(clk), .QN(n5713) );
  EDFD1 \Mem_reg[73][9]  ( .D(n24741), .E(n6404), .CP(clk), .QN(n27075) );
  EDFD1 \Mem_reg[72][9]  ( .D(n24741), .E(n6403), .CP(clk), .QN(n5617) );
  EDFD1 \Mem_reg[71][9]  ( .D(n24741), .E(n6402), .CP(clk), .QN(n5569) );
  EDFD1 \Mem_reg[70][9]  ( .D(n24741), .E(n6401), .CP(clk), .QN(n5521) );
  EDFD1 \Mem_reg[69][9]  ( .D(n24741), .E(n6400), .CP(clk), .QN(n5473) );
  EDFD1 \Mem_reg[68][9]  ( .D(n24741), .E(n6399), .CP(clk), .QN(n5425) );
  EDFD1 \Mem_reg[67][9]  ( .D(n24741), .E(n6398), .CP(clk), .QN(n5377) );
  EDFD1 \Mem_reg[66][9]  ( .D(n24741), .E(n6397), .CP(clk), .QN(n5329) );
  EDFD1 \Mem_reg[65][9]  ( .D(n24741), .E(n6396), .CP(clk), .QN(n15485) );
  EDFD1 \Mem_reg[64][9]  ( .D(n24741), .E(n6395), .CP(clk), .QN(n5233) );
  EDFD1 \Mem_reg[63][9]  ( .D(n24741), .E(n6456), .CP(clk), .QN(n5185) );
  EDFD1 \Mem_reg[62][9]  ( .D(n24741), .E(n6455), .CP(clk), .QN(n5137) );
  EDFD1 \Mem_reg[61][9]  ( .D(n24741), .E(n6454), .CP(clk), .QN(n17954) );
  EDFD1 \Mem_reg[60][9]  ( .D(n24741), .E(n6453), .CP(clk), .QN(n17953) );
  EDFD1 \Mem_reg[59][9]  ( .D(n24741), .E(n6452), .CP(clk), .QN(n4993) );
  EDFD1 \Mem_reg[58][9]  ( .D(n24741), .E(n6451), .CP(clk), .QN(n4945) );
  EDFD1 \Mem_reg[57][9]  ( .D(n24741), .E(n6450), .CP(clk), .QN(n4897) );
  EDFD1 \Mem_reg[56][9]  ( .D(n24741), .E(n6449), .CP(clk), .QN(n4849) );
  EDFD1 \Mem_reg[55][9]  ( .D(n24741), .E(n6448), .CP(clk), .QN(n4801) );
  EDFD1 \Mem_reg[54][9]  ( .D(n24741), .E(n6447), .CP(clk), .QN(n15484) );
  EDFD1 \Mem_reg[53][9]  ( .D(n24741), .E(n6446), .CP(clk), .QN(n4705) );
  EDFD1 \Mem_reg[52][9]  ( .D(n24741), .E(n6445), .CP(clk), .Q(n27072) );
  EDFD1 \Mem_reg[51][9]  ( .D(n24741), .E(n6444), .CP(clk), .QN(n4609) );
  EDFD1 \Mem_reg[50][9]  ( .D(n24741), .E(n6443), .CP(clk), .QN(n4561) );
  EDFD1 \Mem_reg[49][9]  ( .D(n24741), .E(n6442), .CP(clk), .QN(n4513) );
  EDFD1 \Mem_reg[48][9]  ( .D(n24741), .E(n6441), .CP(clk), .QN(n4465) );
  EDFD1 \Mem_reg[47][9]  ( .D(n24741), .E(n6440), .CP(clk), .QN(n4417) );
  EDFD1 \Mem_reg[46][9]  ( .D(n24741), .E(n6439), .CP(clk), .QN(n4369) );
  EDFD1 \Mem_reg[43][9]  ( .D(n24741), .E(n6438), .CP(clk), .QN(n4321) );
  EDFD1 \Mem_reg[42][9]  ( .D(n24741), .E(n6437), .CP(clk), .QN(n4273) );
  EDFD1 \Mem_reg[41][9]  ( .D(n24741), .E(n6436), .CP(clk), .QN(n4225) );
  EDFD1 \Mem_reg[40][9]  ( .D(n24741), .E(n6435), .CP(clk), .QN(n4177) );
  EDFD1 \Mem_reg[39][9]  ( .D(n24741), .E(n6434), .CP(clk), .QN(n4129) );
  EDFD1 \Mem_reg[38][9]  ( .D(n24741), .E(n6433), .CP(clk), .QN(n4081) );
  EDFD1 \Mem_reg[37][9]  ( .D(n24741), .E(n6432), .CP(clk), .QN(n4033) );
  EDFD1 \Mem_reg[36][9]  ( .D(n24741), .E(n6431), .CP(clk), .QN(n3985) );
  EDFD1 \Mem_reg[35][9]  ( .D(n24741), .E(n6430), .CP(clk), .QN(n3937) );
  EDFD1 \Mem_reg[34][9]  ( .D(n24741), .E(n6429), .CP(clk), .QN(n3889) );
  EDFD1 \Mem_reg[33][9]  ( .D(n24741), .E(n6428), .CP(clk), .QN(n3841) );
  EDFD1 \Mem_reg[32][9]  ( .D(n24741), .E(n6427), .CP(clk), .QN(n3793) );
  EDFD1 \Mem_reg[31][9]  ( .D(n24741), .E(n6426), .CP(clk), .QN(n3745) );
  EDFD1 \Mem_reg[30][9]  ( .D(n24741), .E(n6425), .CP(clk), .QN(n3697) );
  EDFD1 \Mem_reg[29][9]  ( .D(n24741), .E(n6424), .CP(clk), .QN(n3649) );
  EDFD1 \Mem_reg[28][9]  ( .D(n24741), .E(n6423), .CP(clk), .QN(n3601) );
  EDFD1 \Mem_reg[27][9]  ( .D(n24741), .E(n6422), .CP(clk), .QN(n3553) );
  EDFD1 \Mem_reg[26][9]  ( .D(n24741), .E(n6421), .CP(clk), .QN(n3505) );
  EDFD1 \Mem_reg[25][9]  ( .D(n24741), .E(n6420), .CP(clk), .QN(n3457) );
  EDFD1 \Mem_reg[24][9]  ( .D(n24741), .E(n6463), .CP(clk), .QN(n3409) );
  EDFD1 \Mem_reg[23][9]  ( .D(n24741), .E(n6464), .CP(clk), .QN(n3361) );
  EDFD1 \Mem_reg[22][9]  ( .D(n24741), .E(n6465), .CP(clk), .QN(n3313) );
  EDFD1 \Mem_reg[21][9]  ( .D(n24741), .E(n6466), .CP(clk), .QN(n3265) );
  EDFD1 \Mem_reg[20][9]  ( .D(n24741), .E(n6467), .CP(clk), .QN(n3217) );
  EDFD1 \Mem_reg[19][9]  ( .D(n24741), .E(n6468), .CP(clk), .QN(n3169) );
  EDFD1 \Mem_reg[18][9]  ( .D(n24741), .E(n6469), .CP(clk), .QN(n3121) );
  EDFD1 \Mem_reg[17][9]  ( .D(n24741), .E(n6470), .CP(clk), .QN(n3073) );
  EDFD1 \Mem_reg[16][9]  ( .D(n24741), .E(n6471), .CP(clk), .QN(n3025) );
  EDFD1 \Mem_reg[15][9]  ( .D(n24741), .E(n6472), .CP(clk), .QN(n2977) );
  EDFD1 \Mem_reg[14][9]  ( .D(n24741), .E(n24720), .CP(clk), .QN(n2929) );
  EDFD1 \Mem_reg[13][9]  ( .D(n24741), .E(n24709), .CP(clk), .QN(n2881) );
  EDFD1 \Mem_reg[12][9]  ( .D(n24741), .E(n24717), .CP(clk), .QN(n2833) );
  EDFD1 \Mem_reg[11][9]  ( .D(n24741), .E(n24707), .CP(clk), .QN(n2785) );
  EDFD1 \Mem_reg[10][9]  ( .D(n24741), .E(n6477), .CP(clk), .QN(n2737) );
  EDFD1 \Mem_reg[9][9]  ( .D(n24741), .E(n24708), .CP(clk), .QN(n2689) );
  EDFD1 \Mem_reg[8][9]  ( .D(n24741), .E(n15642), .CP(clk), .QN(n2641) );
  EDFD1 \Mem_reg[7][9]  ( .D(n24741), .E(n24718), .CP(clk), .QN(n2593) );
  EDFD1 \Mem_reg[6][9]  ( .D(n24741), .E(n24716), .CP(clk), .QN(n2545) );
  EDFD1 \Mem_reg[5][9]  ( .D(n24741), .E(n24719), .CP(clk), .QN(n2497) );
  EDFD1 \Mem_reg[4][9]  ( .D(n24741), .E(n24706), .CP(clk), .QN(n2449) );
  EDFD1 \Mem_reg[3][9]  ( .D(n24741), .E(n24721), .CP(clk), .QN(n2401) );
  EDFD1 \Mem_reg[2][9]  ( .D(n24741), .E(n6460), .CP(clk), .QN(n2353) );
  EDFD1 \Mem_reg[1][9]  ( .D(n24741), .E(n24703), .CP(clk), .QN(n2305) );
  EDFD1 \Mem_reg[0][9]  ( .D(n24741), .E(n24705), .CP(clk), .QN(n2257) );
  EDFD1 \Mem_reg[88][8]  ( .D(n24739), .E(n6419), .CP(clk), .Q(n27069) );
  EDFD1 \Mem_reg[87][8]  ( .D(n24739), .E(n6418), .CP(clk), .QN(n6338) );
  EDFD1 \Mem_reg[86][8]  ( .D(n24739), .E(n6417), .CP(clk), .QN(n24583) );
  EDFD1 \Mem_reg[85][8]  ( .D(n24739), .E(n6416), .CP(clk), .QN(n6242) );
  EDFD1 \Mem_reg[84][8]  ( .D(n24739), .E(n6415), .CP(clk), .QN(n6194) );
  EDFD1 \Mem_reg[83][8]  ( .D(n24739), .E(n6414), .CP(clk), .QN(n6146) );
  EDFD1 \Mem_reg[82][8]  ( .D(n24739), .E(n6413), .CP(clk), .QN(n6098) );
  EDFD1 \Mem_reg[81][8]  ( .D(n24739), .E(n6412), .CP(clk), .QN(n6050) );
  EDFD1 \Mem_reg[80][8]  ( .D(n24739), .E(n6411), .CP(clk), .QN(n6002) );
  EDFD1 \Mem_reg[79][8]  ( .D(n24739), .E(n6410), .CP(clk), .QN(n5954) );
  EDFD1 \Mem_reg[78][8]  ( .D(n24739), .E(n6409), .CP(clk), .QN(n5906) );
  EDFD1 \Mem_reg[77][8]  ( .D(n24739), .E(n6408), .CP(clk), .QN(n5858) );
  EDFD1 \Mem_reg[76][8]  ( .D(n24739), .E(n6407), .CP(clk), .QN(n5810) );
  EDFD1 \Mem_reg[75][8]  ( .D(n24739), .E(n6406), .CP(clk), .QN(n27070) );
  EDFD1 \Mem_reg[74][8]  ( .D(n24739), .E(n6405), .CP(clk), .QN(n5714) );
  EDFD1 \Mem_reg[73][8]  ( .D(n24739), .E(n6404), .CP(clk), .QN(n27071) );
  EDFD1 \Mem_reg[72][8]  ( .D(n24739), .E(n6403), .CP(clk), .QN(n5618) );
  EDFD1 \Mem_reg[71][8]  ( .D(n24739), .E(n6402), .CP(clk), .QN(n5570) );
  EDFD1 \Mem_reg[70][8]  ( .D(n24739), .E(n6401), .CP(clk), .QN(n5522) );
  EDFD1 \Mem_reg[69][8]  ( .D(n24739), .E(n6400), .CP(clk), .QN(n5474) );
  EDFD1 \Mem_reg[68][8]  ( .D(n24739), .E(n6399), .CP(clk), .QN(n5426) );
  EDFD1 \Mem_reg[67][8]  ( .D(n24739), .E(n6398), .CP(clk), .QN(n5378) );
  EDFD1 \Mem_reg[66][8]  ( .D(n24739), .E(n6397), .CP(clk), .QN(n5330) );
  EDFD1 \Mem_reg[65][8]  ( .D(n24739), .E(n6396), .CP(clk), .QN(n15481) );
  EDFD1 \Mem_reg[64][8]  ( .D(n24739), .E(n6395), .CP(clk), .QN(n5234) );
  EDFD1 \Mem_reg[63][8]  ( .D(n24739), .E(n6456), .CP(clk), .QN(n5186) );
  EDFD1 \Mem_reg[62][8]  ( .D(n24739), .E(n6455), .CP(clk), .QN(n5138) );
  EDFD1 \Mem_reg[61][8]  ( .D(n24739), .E(n6454), .CP(clk), .QN(n17951) );
  EDFD1 \Mem_reg[60][8]  ( .D(n24739), .E(n6453), .CP(clk), .QN(n17950) );
  EDFD1 \Mem_reg[59][8]  ( .D(n24739), .E(n6452), .CP(clk), .QN(n4994) );
  EDFD1 \Mem_reg[58][8]  ( .D(n24739), .E(n6451), .CP(clk), .QN(n4946) );
  EDFD1 \Mem_reg[57][8]  ( .D(n24739), .E(n6450), .CP(clk), .QN(n4898) );
  EDFD1 \Mem_reg[56][8]  ( .D(n24739), .E(n6449), .CP(clk), .QN(n4850) );
  EDFD1 \Mem_reg[55][8]  ( .D(n24739), .E(n6448), .CP(clk), .QN(n4802) );
  EDFD1 \Mem_reg[54][8]  ( .D(n24739), .E(n6447), .CP(clk), .QN(n15480) );
  EDFD1 \Mem_reg[53][8]  ( .D(n24739), .E(n6446), .CP(clk), .QN(n4706) );
  EDFD1 \Mem_reg[52][8]  ( .D(n24739), .E(n6445), .CP(clk), .Q(n27068) );
  EDFD1 \Mem_reg[51][8]  ( .D(n24739), .E(n6444), .CP(clk), .QN(n4610) );
  EDFD1 \Mem_reg[50][8]  ( .D(n24739), .E(n6443), .CP(clk), .QN(n4562) );
  EDFD1 \Mem_reg[49][8]  ( .D(n24739), .E(n6442), .CP(clk), .QN(n4514) );
  EDFD1 \Mem_reg[48][8]  ( .D(n24739), .E(n6441), .CP(clk), .QN(n4466) );
  EDFD1 \Mem_reg[47][8]  ( .D(n24739), .E(n6440), .CP(clk), .QN(n4418) );
  EDFD1 \Mem_reg[46][8]  ( .D(n24739), .E(n6439), .CP(clk), .QN(n4370) );
  EDFD1 \Mem_reg[43][8]  ( .D(n24739), .E(n6438), .CP(clk), .QN(n4322) );
  EDFD1 \Mem_reg[42][8]  ( .D(n24739), .E(n6437), .CP(clk), .QN(n4274) );
  EDFD1 \Mem_reg[41][8]  ( .D(n24739), .E(n6436), .CP(clk), .QN(n4226) );
  EDFD1 \Mem_reg[40][8]  ( .D(n24739), .E(n6435), .CP(clk), .QN(n4178) );
  EDFD1 \Mem_reg[39][8]  ( .D(n24739), .E(n6434), .CP(clk), .QN(n4130) );
  EDFD1 \Mem_reg[38][8]  ( .D(n24739), .E(n6433), .CP(clk), .QN(n4082) );
  EDFD1 \Mem_reg[37][8]  ( .D(n24739), .E(n6432), .CP(clk), .QN(n4034) );
  EDFD1 \Mem_reg[36][8]  ( .D(n24739), .E(n6431), .CP(clk), .QN(n3986) );
  EDFD1 \Mem_reg[35][8]  ( .D(n24739), .E(n6430), .CP(clk), .QN(n3938) );
  EDFD1 \Mem_reg[34][8]  ( .D(n24739), .E(n6429), .CP(clk), .QN(n3890) );
  EDFD1 \Mem_reg[33][8]  ( .D(n24739), .E(n6428), .CP(clk), .QN(n3842) );
  EDFD1 \Mem_reg[32][8]  ( .D(n24739), .E(n6427), .CP(clk), .QN(n3794) );
  EDFD1 \Mem_reg[31][8]  ( .D(n24739), .E(n6426), .CP(clk), .QN(n3746) );
  EDFD1 \Mem_reg[30][8]  ( .D(n24739), .E(n6425), .CP(clk), .QN(n3698) );
  EDFD1 \Mem_reg[29][8]  ( .D(n24739), .E(n6424), .CP(clk), .QN(n3650) );
  EDFD1 \Mem_reg[28][8]  ( .D(n24739), .E(n6423), .CP(clk), .QN(n3602) );
  EDFD1 \Mem_reg[27][8]  ( .D(n24739), .E(n6422), .CP(clk), .QN(n3554) );
  EDFD1 \Mem_reg[26][8]  ( .D(n24739), .E(n6421), .CP(clk), .QN(n3506) );
  EDFD1 \Mem_reg[25][8]  ( .D(n24739), .E(n6420), .CP(clk), .QN(n3458) );
  EDFD1 \Mem_reg[24][8]  ( .D(n24739), .E(n6463), .CP(clk), .QN(n3410) );
  EDFD1 \Mem_reg[23][8]  ( .D(n24739), .E(n6464), .CP(clk), .QN(n3362) );
  EDFD1 \Mem_reg[22][8]  ( .D(n24739), .E(n6465), .CP(clk), .QN(n3314) );
  EDFD1 \Mem_reg[21][8]  ( .D(n24739), .E(n6466), .CP(clk), .QN(n3266) );
  EDFD1 \Mem_reg[20][8]  ( .D(n24739), .E(n6467), .CP(clk), .QN(n3218) );
  EDFD1 \Mem_reg[19][8]  ( .D(n24739), .E(n6468), .CP(clk), .QN(n3170) );
  EDFD1 \Mem_reg[18][8]  ( .D(n24739), .E(n6469), .CP(clk), .QN(n3122) );
  EDFD1 \Mem_reg[17][8]  ( .D(n24739), .E(n6470), .CP(clk), .QN(n3074) );
  EDFD1 \Mem_reg[16][8]  ( .D(n24739), .E(n6471), .CP(clk), .QN(n3026) );
  EDFD1 \Mem_reg[15][8]  ( .D(n24739), .E(n6472), .CP(clk), .QN(n2978) );
  EDFD1 \Mem_reg[14][8]  ( .D(n24739), .E(n24720), .CP(clk), .QN(n2930) );
  EDFD1 \Mem_reg[13][8]  ( .D(n24739), .E(n24709), .CP(clk), .QN(n2882) );
  EDFD1 \Mem_reg[12][8]  ( .D(n24739), .E(n24717), .CP(clk), .QN(n2834) );
  EDFD1 \Mem_reg[11][8]  ( .D(n24739), .E(n24707), .CP(clk), .QN(n2786) );
  EDFD1 \Mem_reg[10][8]  ( .D(n24739), .E(n6477), .CP(clk), .QN(n2738) );
  EDFD1 \Mem_reg[9][8]  ( .D(n24739), .E(n24708), .CP(clk), .QN(n2690) );
  EDFD1 \Mem_reg[8][8]  ( .D(n24739), .E(n15642), .CP(clk), .QN(n2642) );
  EDFD1 \Mem_reg[7][8]  ( .D(n24739), .E(n24718), .CP(clk), .QN(n2594) );
  EDFD1 \Mem_reg[6][8]  ( .D(n24739), .E(n24716), .CP(clk), .QN(n2546) );
  EDFD1 \Mem_reg[5][8]  ( .D(n24739), .E(n24719), .CP(clk), .QN(n2498) );
  EDFD1 \Mem_reg[4][8]  ( .D(n24739), .E(n24706), .CP(clk), .QN(n2450) );
  EDFD1 \Mem_reg[3][8]  ( .D(n24739), .E(n24721), .CP(clk), .QN(n2402) );
  EDFD1 \Mem_reg[2][8]  ( .D(n24739), .E(n6460), .CP(clk), .QN(n2354) );
  EDFD1 \Mem_reg[1][8]  ( .D(n24739), .E(n24703), .CP(clk), .QN(n2306) );
  EDFD1 \Mem_reg[0][8]  ( .D(n24739), .E(n24705), .CP(clk), .QN(n2258) );
  EDFD1 \Mem_reg[88][7]  ( .D(n24737), .E(n6419), .CP(clk), .Q(n27065) );
  EDFD1 \Mem_reg[87][7]  ( .D(n24737), .E(n6418), .CP(clk), .QN(n6339) );
  EDFD1 \Mem_reg[86][7]  ( .D(n24737), .E(n6417), .CP(clk), .QN(n24580) );
  EDFD1 \Mem_reg[85][7]  ( .D(n24737), .E(n6416), .CP(clk), .QN(n6243) );
  EDFD1 \Mem_reg[84][7]  ( .D(n24737), .E(n6415), .CP(clk), .QN(n6195) );
  EDFD1 \Mem_reg[83][7]  ( .D(n24737), .E(n6414), .CP(clk), .QN(n6147) );
  EDFD1 \Mem_reg[82][7]  ( .D(n24737), .E(n6413), .CP(clk), .QN(n6099) );
  EDFD1 \Mem_reg[81][7]  ( .D(n24737), .E(n6412), .CP(clk), .QN(n6051) );
  EDFD1 \Mem_reg[80][7]  ( .D(n24737), .E(n6411), .CP(clk), .QN(n6003) );
  EDFD1 \Mem_reg[79][7]  ( .D(n24737), .E(n6410), .CP(clk), .QN(n5955) );
  EDFD1 \Mem_reg[78][7]  ( .D(n24737), .E(n6409), .CP(clk), .QN(n5907) );
  EDFD1 \Mem_reg[77][7]  ( .D(n24737), .E(n6408), .CP(clk), .QN(n5859) );
  EDFD1 \Mem_reg[76][7]  ( .D(n24737), .E(n6407), .CP(clk), .QN(n5811) );
  EDFD1 \Mem_reg[75][7]  ( .D(n24737), .E(n6406), .CP(clk), .QN(n27066) );
  EDFD1 \Mem_reg[74][7]  ( .D(n24737), .E(n6405), .CP(clk), .QN(n5715) );
  EDFD1 \Mem_reg[73][7]  ( .D(n24737), .E(n6404), .CP(clk), .QN(n27067) );
  EDFD1 \Mem_reg[72][7]  ( .D(n24737), .E(n6403), .CP(clk), .QN(n5619) );
  EDFD1 \Mem_reg[71][7]  ( .D(n24737), .E(n6402), .CP(clk), .QN(n5571) );
  EDFD1 \Mem_reg[70][7]  ( .D(n24737), .E(n6401), .CP(clk), .QN(n5523) );
  EDFD1 \Mem_reg[69][7]  ( .D(n24737), .E(n6400), .CP(clk), .QN(n5475) );
  EDFD1 \Mem_reg[68][7]  ( .D(n24737), .E(n6399), .CP(clk), .QN(n5427) );
  EDFD1 \Mem_reg[67][7]  ( .D(n24737), .E(n6398), .CP(clk), .QN(n5379) );
  EDFD1 \Mem_reg[66][7]  ( .D(n24737), .E(n6397), .CP(clk), .QN(n5331) );
  EDFD1 \Mem_reg[65][7]  ( .D(n24737), .E(n6396), .CP(clk), .QN(n15477) );
  EDFD1 \Mem_reg[64][7]  ( .D(n24737), .E(n6395), .CP(clk), .QN(n5235) );
  EDFD1 \Mem_reg[63][7]  ( .D(n24737), .E(n6456), .CP(clk), .QN(n5187) );
  EDFD1 \Mem_reg[62][7]  ( .D(n24737), .E(n6455), .CP(clk), .QN(n5139) );
  EDFD1 \Mem_reg[61][7]  ( .D(n24737), .E(n6454), .CP(clk), .QN(n17948) );
  EDFD1 \Mem_reg[60][7]  ( .D(n24737), .E(n6453), .CP(clk), .QN(n17947) );
  EDFD1 \Mem_reg[59][7]  ( .D(n24737), .E(n6452), .CP(clk), .QN(n4995) );
  EDFD1 \Mem_reg[58][7]  ( .D(n24737), .E(n6451), .CP(clk), .QN(n4947) );
  EDFD1 \Mem_reg[57][7]  ( .D(n24737), .E(n6450), .CP(clk), .QN(n4899) );
  EDFD1 \Mem_reg[56][7]  ( .D(n24737), .E(n6449), .CP(clk), .QN(n4851) );
  EDFD1 \Mem_reg[55][7]  ( .D(n24737), .E(n6448), .CP(clk), .QN(n4803) );
  EDFD1 \Mem_reg[54][7]  ( .D(n24737), .E(n6447), .CP(clk), .QN(n15476) );
  EDFD1 \Mem_reg[53][7]  ( .D(n24737), .E(n6446), .CP(clk), .QN(n4707) );
  EDFD1 \Mem_reg[52][7]  ( .D(n24737), .E(n6445), .CP(clk), .Q(n27064) );
  EDFD1 \Mem_reg[51][7]  ( .D(n24737), .E(n6444), .CP(clk), .QN(n4611) );
  EDFD1 \Mem_reg[50][7]  ( .D(n24737), .E(n6443), .CP(clk), .QN(n4563) );
  EDFD1 \Mem_reg[49][7]  ( .D(n24737), .E(n6442), .CP(clk), .QN(n4515) );
  EDFD1 \Mem_reg[48][7]  ( .D(n24737), .E(n6441), .CP(clk), .QN(n4467) );
  EDFD1 \Mem_reg[47][7]  ( .D(n24737), .E(n6440), .CP(clk), .QN(n4419) );
  EDFD1 \Mem_reg[46][7]  ( .D(n24737), .E(n6439), .CP(clk), .QN(n4371) );
  EDFD1 \Mem_reg[43][7]  ( .D(n24737), .E(n6438), .CP(clk), .QN(n4323) );
  EDFD1 \Mem_reg[42][7]  ( .D(n24737), .E(n6437), .CP(clk), .QN(n4275) );
  EDFD1 \Mem_reg[41][7]  ( .D(n24737), .E(n6436), .CP(clk), .QN(n4227) );
  EDFD1 \Mem_reg[40][7]  ( .D(n24737), .E(n6435), .CP(clk), .QN(n4179) );
  EDFD1 \Mem_reg[39][7]  ( .D(n24737), .E(n6434), .CP(clk), .QN(n4131) );
  EDFD1 \Mem_reg[38][7]  ( .D(n24737), .E(n6433), .CP(clk), .QN(n4083) );
  EDFD1 \Mem_reg[37][7]  ( .D(n24737), .E(n6432), .CP(clk), .QN(n4035) );
  EDFD1 \Mem_reg[36][7]  ( .D(n24737), .E(n6431), .CP(clk), .QN(n3987) );
  EDFD1 \Mem_reg[35][7]  ( .D(n24737), .E(n6430), .CP(clk), .QN(n3939) );
  EDFD1 \Mem_reg[34][7]  ( .D(n24737), .E(n6429), .CP(clk), .QN(n3891) );
  EDFD1 \Mem_reg[33][7]  ( .D(n24737), .E(n6428), .CP(clk), .QN(n3843) );
  EDFD1 \Mem_reg[32][7]  ( .D(n24737), .E(n6427), .CP(clk), .QN(n3795) );
  EDFD1 \Mem_reg[31][7]  ( .D(n24737), .E(n6426), .CP(clk), .QN(n3747) );
  EDFD1 \Mem_reg[30][7]  ( .D(n24737), .E(n6425), .CP(clk), .QN(n3699) );
  EDFD1 \Mem_reg[29][7]  ( .D(n24737), .E(n6424), .CP(clk), .QN(n3651) );
  EDFD1 \Mem_reg[28][7]  ( .D(n24737), .E(n6423), .CP(clk), .QN(n3603) );
  EDFD1 \Mem_reg[27][7]  ( .D(n24737), .E(n6422), .CP(clk), .QN(n3555) );
  EDFD1 \Mem_reg[26][7]  ( .D(n24737), .E(n6421), .CP(clk), .QN(n3507) );
  EDFD1 \Mem_reg[25][7]  ( .D(n24737), .E(n6420), .CP(clk), .QN(n3459) );
  EDFD1 \Mem_reg[24][7]  ( .D(n24737), .E(n6463), .CP(clk), .QN(n3411) );
  EDFD1 \Mem_reg[23][7]  ( .D(n24737), .E(n6464), .CP(clk), .QN(n3363) );
  EDFD1 \Mem_reg[22][7]  ( .D(n24737), .E(n6465), .CP(clk), .QN(n3315) );
  EDFD1 \Mem_reg[21][7]  ( .D(n24737), .E(n6466), .CP(clk), .QN(n3267) );
  EDFD1 \Mem_reg[20][7]  ( .D(n24737), .E(n6467), .CP(clk), .QN(n3219) );
  EDFD1 \Mem_reg[19][7]  ( .D(n24737), .E(n6468), .CP(clk), .QN(n3171) );
  EDFD1 \Mem_reg[18][7]  ( .D(n24737), .E(n6469), .CP(clk), .QN(n3123) );
  EDFD1 \Mem_reg[17][7]  ( .D(n24737), .E(n6470), .CP(clk), .QN(n3075) );
  EDFD1 \Mem_reg[16][7]  ( .D(n24737), .E(n6471), .CP(clk), .QN(n3027) );
  EDFD1 \Mem_reg[15][7]  ( .D(n24737), .E(n6472), .CP(clk), .QN(n2979) );
  EDFD1 \Mem_reg[14][7]  ( .D(n24737), .E(n24720), .CP(clk), .QN(n2931) );
  EDFD1 \Mem_reg[13][7]  ( .D(n24737), .E(n24709), .CP(clk), .QN(n2883) );
  EDFD1 \Mem_reg[12][7]  ( .D(n24737), .E(n24717), .CP(clk), .QN(n2835) );
  EDFD1 \Mem_reg[11][7]  ( .D(n24737), .E(n24707), .CP(clk), .QN(n2787) );
  EDFD1 \Mem_reg[10][7]  ( .D(n24737), .E(n6477), .CP(clk), .QN(n2739) );
  EDFD1 \Mem_reg[9][7]  ( .D(n24737), .E(n24708), .CP(clk), .QN(n2691) );
  EDFD1 \Mem_reg[8][7]  ( .D(n24737), .E(n15642), .CP(clk), .QN(n2643) );
  EDFD1 \Mem_reg[7][7]  ( .D(n24737), .E(n24718), .CP(clk), .QN(n2595) );
  EDFD1 \Mem_reg[6][7]  ( .D(n24737), .E(n24716), .CP(clk), .QN(n2547) );
  EDFD1 \Mem_reg[5][7]  ( .D(n24737), .E(n24719), .CP(clk), .QN(n2499) );
  EDFD1 \Mem_reg[4][7]  ( .D(n24737), .E(n24706), .CP(clk), .QN(n2451) );
  EDFD1 \Mem_reg[3][7]  ( .D(n24737), .E(n24721), .CP(clk), .QN(n2403) );
  EDFD1 \Mem_reg[2][7]  ( .D(n24737), .E(n6460), .CP(clk), .QN(n2355) );
  EDFD1 \Mem_reg[1][7]  ( .D(n24737), .E(n24703), .CP(clk), .QN(n2307) );
  EDFD1 \Mem_reg[0][7]  ( .D(n24737), .E(n24705), .CP(clk), .QN(n2259) );
  EDFD1 \Mem_reg[88][6]  ( .D(n24735), .E(n6419), .CP(clk), .Q(n27061) );
  EDFD1 \Mem_reg[87][6]  ( .D(n24735), .E(n6418), .CP(clk), .QN(n6340) );
  EDFD1 \Mem_reg[86][6]  ( .D(n24735), .E(n6417), .CP(clk), .QN(n24577) );
  EDFD1 \Mem_reg[85][6]  ( .D(n24735), .E(n6416), .CP(clk), .QN(n6244) );
  EDFD1 \Mem_reg[84][6]  ( .D(n24735), .E(n6415), .CP(clk), .QN(n6196) );
  EDFD1 \Mem_reg[83][6]  ( .D(n24735), .E(n6414), .CP(clk), .QN(n6148) );
  EDFD1 \Mem_reg[82][6]  ( .D(n24735), .E(n6413), .CP(clk), .QN(n6100) );
  EDFD1 \Mem_reg[81][6]  ( .D(n24735), .E(n6412), .CP(clk), .QN(n6052) );
  EDFD1 \Mem_reg[80][6]  ( .D(n24735), .E(n6411), .CP(clk), .QN(n6004) );
  EDFD1 \Mem_reg[79][6]  ( .D(n24735), .E(n6410), .CP(clk), .QN(n5956) );
  EDFD1 \Mem_reg[78][6]  ( .D(n24735), .E(n6409), .CP(clk), .QN(n5908) );
  EDFD1 \Mem_reg[77][6]  ( .D(n24735), .E(n6408), .CP(clk), .QN(n5860) );
  EDFD1 \Mem_reg[76][6]  ( .D(n24735), .E(n6407), .CP(clk), .QN(n5812) );
  EDFD1 \Mem_reg[75][6]  ( .D(n24735), .E(n6406), .CP(clk), .QN(n27062) );
  EDFD1 \Mem_reg[74][6]  ( .D(n24735), .E(n6405), .CP(clk), .QN(n5716) );
  EDFD1 \Mem_reg[73][6]  ( .D(n24735), .E(n6404), .CP(clk), .QN(n27063) );
  EDFD1 \Mem_reg[72][6]  ( .D(n24735), .E(n6403), .CP(clk), .QN(n5620) );
  EDFD1 \Mem_reg[71][6]  ( .D(n24735), .E(n6402), .CP(clk), .QN(n5572) );
  EDFD1 \Mem_reg[70][6]  ( .D(n24735), .E(n6401), .CP(clk), .QN(n5524) );
  EDFD1 \Mem_reg[69][6]  ( .D(n24735), .E(n6400), .CP(clk), .QN(n5476) );
  EDFD1 \Mem_reg[68][6]  ( .D(n24735), .E(n6399), .CP(clk), .QN(n5428) );
  EDFD1 \Mem_reg[67][6]  ( .D(n24735), .E(n6398), .CP(clk), .QN(n5380) );
  EDFD1 \Mem_reg[66][6]  ( .D(n24735), .E(n6397), .CP(clk), .QN(n5332) );
  EDFD1 \Mem_reg[65][6]  ( .D(n24735), .E(n6396), .CP(clk), .QN(n15473) );
  EDFD1 \Mem_reg[64][6]  ( .D(n24735), .E(n6395), .CP(clk), .QN(n5236) );
  EDFD1 \Mem_reg[63][6]  ( .D(n24735), .E(n6456), .CP(clk), .QN(n5188) );
  EDFD1 \Mem_reg[62][6]  ( .D(n24735), .E(n6455), .CP(clk), .QN(n5140) );
  EDFD1 \Mem_reg[61][6]  ( .D(n24735), .E(n6454), .CP(clk), .QN(n17945) );
  EDFD1 \Mem_reg[60][6]  ( .D(n24735), .E(n6453), .CP(clk), .QN(n17944) );
  EDFD1 \Mem_reg[59][6]  ( .D(n24735), .E(n6452), .CP(clk), .QN(n4996) );
  EDFD1 \Mem_reg[58][6]  ( .D(n24735), .E(n6451), .CP(clk), .QN(n4948) );
  EDFD1 \Mem_reg[57][6]  ( .D(n24735), .E(n6450), .CP(clk), .QN(n4900) );
  EDFD1 \Mem_reg[56][6]  ( .D(n24735), .E(n6449), .CP(clk), .QN(n4852) );
  EDFD1 \Mem_reg[55][6]  ( .D(n24735), .E(n6448), .CP(clk), .QN(n4804) );
  EDFD1 \Mem_reg[54][6]  ( .D(n24735), .E(n6447), .CP(clk), .QN(n15472) );
  EDFD1 \Mem_reg[53][6]  ( .D(n24735), .E(n6446), .CP(clk), .QN(n4708) );
  EDFD1 \Mem_reg[52][6]  ( .D(n24735), .E(n6445), .CP(clk), .Q(n27060) );
  EDFD1 \Mem_reg[51][6]  ( .D(n24735), .E(n6444), .CP(clk), .QN(n4612) );
  EDFD1 \Mem_reg[50][6]  ( .D(n24735), .E(n6443), .CP(clk), .QN(n4564) );
  EDFD1 \Mem_reg[49][6]  ( .D(n24735), .E(n6442), .CP(clk), .QN(n4516) );
  EDFD1 \Mem_reg[48][6]  ( .D(n24735), .E(n6441), .CP(clk), .QN(n4468) );
  EDFD1 \Mem_reg[47][6]  ( .D(n24735), .E(n6440), .CP(clk), .QN(n4420) );
  EDFD1 \Mem_reg[46][6]  ( .D(n24735), .E(n6439), .CP(clk), .QN(n4372) );
  EDFD1 \Mem_reg[43][6]  ( .D(n24735), .E(n6438), .CP(clk), .QN(n4324) );
  EDFD1 \Mem_reg[42][6]  ( .D(n24735), .E(n6437), .CP(clk), .QN(n4276) );
  EDFD1 \Mem_reg[41][6]  ( .D(n24735), .E(n6436), .CP(clk), .QN(n4228) );
  EDFD1 \Mem_reg[40][6]  ( .D(n24735), .E(n6435), .CP(clk), .QN(n4180) );
  EDFD1 \Mem_reg[39][6]  ( .D(n24735), .E(n6434), .CP(clk), .QN(n4132) );
  EDFD1 \Mem_reg[38][6]  ( .D(n24735), .E(n6433), .CP(clk), .QN(n4084) );
  EDFD1 \Mem_reg[37][6]  ( .D(n24735), .E(n6432), .CP(clk), .QN(n4036) );
  EDFD1 \Mem_reg[36][6]  ( .D(n24735), .E(n6431), .CP(clk), .QN(n3988) );
  EDFD1 \Mem_reg[35][6]  ( .D(n24735), .E(n6430), .CP(clk), .QN(n3940) );
  EDFD1 \Mem_reg[34][6]  ( .D(n24735), .E(n6429), .CP(clk), .QN(n3892) );
  EDFD1 \Mem_reg[33][6]  ( .D(n24735), .E(n6428), .CP(clk), .QN(n3844) );
  EDFD1 \Mem_reg[32][6]  ( .D(n24735), .E(n6427), .CP(clk), .QN(n3796) );
  EDFD1 \Mem_reg[31][6]  ( .D(n24735), .E(n6426), .CP(clk), .QN(n3748) );
  EDFD1 \Mem_reg[30][6]  ( .D(n24735), .E(n6425), .CP(clk), .QN(n3700) );
  EDFD1 \Mem_reg[29][6]  ( .D(n24735), .E(n6424), .CP(clk), .QN(n3652) );
  EDFD1 \Mem_reg[28][6]  ( .D(n24735), .E(n6423), .CP(clk), .QN(n3604) );
  EDFD1 \Mem_reg[27][6]  ( .D(n24735), .E(n6422), .CP(clk), .QN(n3556) );
  EDFD1 \Mem_reg[26][6]  ( .D(n24735), .E(n6421), .CP(clk), .QN(n3508) );
  EDFD1 \Mem_reg[25][6]  ( .D(n24735), .E(n6420), .CP(clk), .QN(n3460) );
  EDFD1 \Mem_reg[24][6]  ( .D(n24735), .E(n6463), .CP(clk), .QN(n3412) );
  EDFD1 \Mem_reg[23][6]  ( .D(n24735), .E(n6464), .CP(clk), .QN(n3364) );
  EDFD1 \Mem_reg[22][6]  ( .D(n24735), .E(n6465), .CP(clk), .QN(n3316) );
  EDFD1 \Mem_reg[21][6]  ( .D(n24735), .E(n6466), .CP(clk), .QN(n3268) );
  EDFD1 \Mem_reg[20][6]  ( .D(n24735), .E(n6467), .CP(clk), .QN(n3220) );
  EDFD1 \Mem_reg[19][6]  ( .D(n24735), .E(n6468), .CP(clk), .QN(n3172) );
  EDFD1 \Mem_reg[18][6]  ( .D(n24735), .E(n6469), .CP(clk), .QN(n3124) );
  EDFD1 \Mem_reg[17][6]  ( .D(n24735), .E(n6470), .CP(clk), .QN(n3076) );
  EDFD1 \Mem_reg[16][6]  ( .D(n24735), .E(n6471), .CP(clk), .QN(n3028) );
  EDFD1 \Mem_reg[15][6]  ( .D(n24735), .E(n6472), .CP(clk), .QN(n2980) );
  EDFD1 \Mem_reg[14][6]  ( .D(n24735), .E(n24720), .CP(clk), .QN(n2932) );
  EDFD1 \Mem_reg[13][6]  ( .D(n24735), .E(n24709), .CP(clk), .QN(n2884) );
  EDFD1 \Mem_reg[12][6]  ( .D(n24735), .E(n24717), .CP(clk), .QN(n2836) );
  EDFD1 \Mem_reg[11][6]  ( .D(n24735), .E(n24707), .CP(clk), .QN(n2788) );
  EDFD1 \Mem_reg[10][6]  ( .D(n24735), .E(n6477), .CP(clk), .QN(n2740) );
  EDFD1 \Mem_reg[9][6]  ( .D(n24735), .E(n24708), .CP(clk), .QN(n2692) );
  EDFD1 \Mem_reg[8][6]  ( .D(n24735), .E(n15642), .CP(clk), .QN(n2644) );
  EDFD1 \Mem_reg[7][6]  ( .D(n24735), .E(n24718), .CP(clk), .QN(n2596) );
  EDFD1 \Mem_reg[6][6]  ( .D(n24735), .E(n24716), .CP(clk), .QN(n2548) );
  EDFD1 \Mem_reg[5][6]  ( .D(n24735), .E(n24719), .CP(clk), .QN(n2500) );
  EDFD1 \Mem_reg[4][6]  ( .D(n24735), .E(n24706), .CP(clk), .QN(n2452) );
  EDFD1 \Mem_reg[3][6]  ( .D(n24735), .E(n24721), .CP(clk), .QN(n2404) );
  EDFD1 \Mem_reg[2][6]  ( .D(n24735), .E(n6460), .CP(clk), .QN(n2356) );
  EDFD1 \Mem_reg[1][6]  ( .D(n24735), .E(n24703), .CP(clk), .QN(n2308) );
  EDFD1 \Mem_reg[0][6]  ( .D(n24735), .E(n24705), .CP(clk), .QN(n2260) );
  EDFD1 \Mem_reg[88][5]  ( .D(n24733), .E(n6419), .CP(clk), .Q(n27057) );
  EDFD1 \Mem_reg[87][5]  ( .D(n24733), .E(n6418), .CP(clk), .QN(n6341) );
  EDFD1 \Mem_reg[86][5]  ( .D(n24733), .E(n6417), .CP(clk), .QN(n24574) );
  EDFD1 \Mem_reg[85][5]  ( .D(n24733), .E(n6416), .CP(clk), .QN(n6245) );
  EDFD1 \Mem_reg[84][5]  ( .D(n24733), .E(n6415), .CP(clk), .QN(n6197) );
  EDFD1 \Mem_reg[83][5]  ( .D(n24733), .E(n6414), .CP(clk), .QN(n6149) );
  EDFD1 \Mem_reg[82][5]  ( .D(n24733), .E(n6413), .CP(clk), .QN(n6101) );
  EDFD1 \Mem_reg[81][5]  ( .D(n24733), .E(n6412), .CP(clk), .QN(n6053) );
  EDFD1 \Mem_reg[80][5]  ( .D(n24733), .E(n6411), .CP(clk), .QN(n6005) );
  EDFD1 \Mem_reg[79][5]  ( .D(n24733), .E(n6410), .CP(clk), .QN(n5957) );
  EDFD1 \Mem_reg[78][5]  ( .D(n24733), .E(n6409), .CP(clk), .QN(n5909) );
  EDFD1 \Mem_reg[77][5]  ( .D(n24733), .E(n6408), .CP(clk), .QN(n5861) );
  EDFD1 \Mem_reg[76][5]  ( .D(n24733), .E(n6407), .CP(clk), .QN(n5813) );
  EDFD1 \Mem_reg[75][5]  ( .D(n24733), .E(n6406), .CP(clk), .QN(n27058) );
  EDFD1 \Mem_reg[74][5]  ( .D(n24733), .E(n6405), .CP(clk), .QN(n5717) );
  EDFD1 \Mem_reg[73][5]  ( .D(n24733), .E(n6404), .CP(clk), .QN(n27059) );
  EDFD1 \Mem_reg[72][5]  ( .D(n24733), .E(n6403), .CP(clk), .QN(n5621) );
  EDFD1 \Mem_reg[71][5]  ( .D(n24733), .E(n6402), .CP(clk), .QN(n5573) );
  EDFD1 \Mem_reg[70][5]  ( .D(n24733), .E(n6401), .CP(clk), .QN(n5525) );
  EDFD1 \Mem_reg[69][5]  ( .D(n24733), .E(n6400), .CP(clk), .QN(n5477) );
  EDFD1 \Mem_reg[68][5]  ( .D(n24733), .E(n6399), .CP(clk), .QN(n5429) );
  EDFD1 \Mem_reg[67][5]  ( .D(n24733), .E(n6398), .CP(clk), .QN(n5381) );
  EDFD1 \Mem_reg[66][5]  ( .D(n24733), .E(n6397), .CP(clk), .QN(n5333) );
  EDFD1 \Mem_reg[65][5]  ( .D(n24733), .E(n6396), .CP(clk), .QN(n15469) );
  EDFD1 \Mem_reg[64][5]  ( .D(n24733), .E(n6395), .CP(clk), .QN(n5237) );
  EDFD1 \Mem_reg[63][5]  ( .D(n24733), .E(n6456), .CP(clk), .QN(n5189) );
  EDFD1 \Mem_reg[62][5]  ( .D(n24733), .E(n6455), .CP(clk), .QN(n5141) );
  EDFD1 \Mem_reg[61][5]  ( .D(n24733), .E(n6454), .CP(clk), .QN(n17942) );
  EDFD1 \Mem_reg[60][5]  ( .D(n24733), .E(n6453), .CP(clk), .QN(n17941) );
  EDFD1 \Mem_reg[59][5]  ( .D(n24733), .E(n6452), .CP(clk), .QN(n4997) );
  EDFD1 \Mem_reg[58][5]  ( .D(n24733), .E(n6451), .CP(clk), .QN(n4949) );
  EDFD1 \Mem_reg[57][5]  ( .D(n24733), .E(n6450), .CP(clk), .QN(n4901) );
  EDFD1 \Mem_reg[56][5]  ( .D(n24733), .E(n6449), .CP(clk), .QN(n4853) );
  EDFD1 \Mem_reg[55][5]  ( .D(n24733), .E(n6448), .CP(clk), .QN(n4805) );
  EDFD1 \Mem_reg[54][5]  ( .D(n24733), .E(n6447), .CP(clk), .QN(n15468) );
  EDFD1 \Mem_reg[53][5]  ( .D(n24733), .E(n6446), .CP(clk), .QN(n4709) );
  EDFD1 \Mem_reg[52][5]  ( .D(n24733), .E(n6445), .CP(clk), .Q(n27056) );
  EDFD1 \Mem_reg[51][5]  ( .D(n24733), .E(n6444), .CP(clk), .QN(n4613) );
  EDFD1 \Mem_reg[50][5]  ( .D(n24733), .E(n6443), .CP(clk), .QN(n4565) );
  EDFD1 \Mem_reg[49][5]  ( .D(n24733), .E(n6442), .CP(clk), .QN(n4517) );
  EDFD1 \Mem_reg[48][5]  ( .D(n24733), .E(n6441), .CP(clk), .QN(n4469) );
  EDFD1 \Mem_reg[47][5]  ( .D(n24733), .E(n6440), .CP(clk), .QN(n4421) );
  EDFD1 \Mem_reg[46][5]  ( .D(n24733), .E(n6439), .CP(clk), .QN(n4373) );
  EDFD1 \Mem_reg[43][5]  ( .D(n24733), .E(n6438), .CP(clk), .QN(n4325) );
  EDFD1 \Mem_reg[42][5]  ( .D(n24733), .E(n6437), .CP(clk), .QN(n4277) );
  EDFD1 \Mem_reg[41][5]  ( .D(n24733), .E(n6436), .CP(clk), .QN(n4229) );
  EDFD1 \Mem_reg[40][5]  ( .D(n24733), .E(n6435), .CP(clk), .QN(n4181) );
  EDFD1 \Mem_reg[39][5]  ( .D(n24733), .E(n6434), .CP(clk), .QN(n4133) );
  EDFD1 \Mem_reg[38][5]  ( .D(n24733), .E(n6433), .CP(clk), .QN(n4085) );
  EDFD1 \Mem_reg[37][5]  ( .D(n24733), .E(n6432), .CP(clk), .QN(n4037) );
  EDFD1 \Mem_reg[36][5]  ( .D(n24733), .E(n6431), .CP(clk), .QN(n3989) );
  EDFD1 \Mem_reg[35][5]  ( .D(n24733), .E(n6430), .CP(clk), .QN(n3941) );
  EDFD1 \Mem_reg[34][5]  ( .D(n24733), .E(n6429), .CP(clk), .QN(n3893) );
  EDFD1 \Mem_reg[33][5]  ( .D(n24733), .E(n6428), .CP(clk), .QN(n3845) );
  EDFD1 \Mem_reg[32][5]  ( .D(n24733), .E(n6427), .CP(clk), .QN(n3797) );
  EDFD1 \Mem_reg[31][5]  ( .D(n24733), .E(n6426), .CP(clk), .QN(n3749) );
  EDFD1 \Mem_reg[30][5]  ( .D(n24733), .E(n6425), .CP(clk), .QN(n3701) );
  EDFD1 \Mem_reg[29][5]  ( .D(n24733), .E(n6424), .CP(clk), .QN(n3653) );
  EDFD1 \Mem_reg[28][5]  ( .D(n24733), .E(n6423), .CP(clk), .QN(n3605) );
  EDFD1 \Mem_reg[27][5]  ( .D(n24733), .E(n6422), .CP(clk), .QN(n3557) );
  EDFD1 \Mem_reg[26][5]  ( .D(n24733), .E(n6421), .CP(clk), .QN(n3509) );
  EDFD1 \Mem_reg[25][5]  ( .D(n24733), .E(n6420), .CP(clk), .QN(n3461) );
  EDFD1 \Mem_reg[24][5]  ( .D(n24733), .E(n6463), .CP(clk), .QN(n3413) );
  EDFD1 \Mem_reg[23][5]  ( .D(n24733), .E(n6464), .CP(clk), .QN(n3365) );
  EDFD1 \Mem_reg[22][5]  ( .D(n24733), .E(n6465), .CP(clk), .QN(n3317) );
  EDFD1 \Mem_reg[21][5]  ( .D(n24733), .E(n6466), .CP(clk), .QN(n3269) );
  EDFD1 \Mem_reg[20][5]  ( .D(n24733), .E(n6467), .CP(clk), .QN(n3221) );
  EDFD1 \Mem_reg[19][5]  ( .D(n24733), .E(n6468), .CP(clk), .QN(n3173) );
  EDFD1 \Mem_reg[18][5]  ( .D(n24733), .E(n6469), .CP(clk), .QN(n3125) );
  EDFD1 \Mem_reg[17][5]  ( .D(n24733), .E(n6470), .CP(clk), .QN(n3077) );
  EDFD1 \Mem_reg[16][5]  ( .D(n24733), .E(n6471), .CP(clk), .QN(n3029) );
  EDFD1 \Mem_reg[15][5]  ( .D(n24733), .E(n6472), .CP(clk), .QN(n2981) );
  EDFD1 \Mem_reg[14][5]  ( .D(n24733), .E(n24720), .CP(clk), .QN(n2933) );
  EDFD1 \Mem_reg[13][5]  ( .D(n24733), .E(n24709), .CP(clk), .QN(n2885) );
  EDFD1 \Mem_reg[12][5]  ( .D(n24733), .E(n24717), .CP(clk), .QN(n2837) );
  EDFD1 \Mem_reg[11][5]  ( .D(n24733), .E(n24707), .CP(clk), .QN(n2789) );
  EDFD1 \Mem_reg[10][5]  ( .D(n24733), .E(n6477), .CP(clk), .QN(n2741) );
  EDFD1 \Mem_reg[9][5]  ( .D(n24733), .E(n24708), .CP(clk), .QN(n2693) );
  EDFD1 \Mem_reg[8][5]  ( .D(n24733), .E(n15642), .CP(clk), .QN(n2645) );
  EDFD1 \Mem_reg[7][5]  ( .D(n24733), .E(n24718), .CP(clk), .QN(n2597) );
  EDFD1 \Mem_reg[6][5]  ( .D(n24733), .E(n24716), .CP(clk), .QN(n2549) );
  EDFD1 \Mem_reg[5][5]  ( .D(n24733), .E(n24719), .CP(clk), .QN(n2501) );
  EDFD1 \Mem_reg[4][5]  ( .D(n24733), .E(n24706), .CP(clk), .QN(n2453) );
  EDFD1 \Mem_reg[3][5]  ( .D(n24733), .E(n24721), .CP(clk), .QN(n2405) );
  EDFD1 \Mem_reg[2][5]  ( .D(n24733), .E(n6460), .CP(clk), .QN(n2357) );
  EDFD1 \Mem_reg[1][5]  ( .D(n24733), .E(n24703), .CP(clk), .QN(n2309) );
  EDFD1 \Mem_reg[0][5]  ( .D(n24733), .E(n24705), .CP(clk), .QN(n2261) );
  EDFD1 \Mem_reg[88][4]  ( .D(n24731), .E(n6419), .CP(clk), .Q(n27053) );
  EDFD1 \Mem_reg[87][4]  ( .D(n24731), .E(n6418), .CP(clk), .QN(n6342) );
  EDFD1 \Mem_reg[86][4]  ( .D(n24731), .E(n6417), .CP(clk), .QN(n24571) );
  EDFD1 \Mem_reg[85][4]  ( .D(n24731), .E(n6416), .CP(clk), .QN(n6246) );
  EDFD1 \Mem_reg[84][4]  ( .D(n24731), .E(n6415), .CP(clk), .QN(n6198) );
  EDFD1 \Mem_reg[83][4]  ( .D(n24731), .E(n6414), .CP(clk), .QN(n6150) );
  EDFD1 \Mem_reg[82][4]  ( .D(n24731), .E(n6413), .CP(clk), .QN(n6102) );
  EDFD1 \Mem_reg[81][4]  ( .D(n24731), .E(n6412), .CP(clk), .QN(n6054) );
  EDFD1 \Mem_reg[80][4]  ( .D(n24731), .E(n6411), .CP(clk), .QN(n6006) );
  EDFD1 \Mem_reg[79][4]  ( .D(n24731), .E(n6410), .CP(clk), .QN(n5958) );
  EDFD1 \Mem_reg[78][4]  ( .D(n24731), .E(n6409), .CP(clk), .QN(n5910) );
  EDFD1 \Mem_reg[77][4]  ( .D(n24731), .E(n6408), .CP(clk), .QN(n5862) );
  EDFD1 \Mem_reg[76][4]  ( .D(n24731), .E(n6407), .CP(clk), .QN(n5814) );
  EDFD1 \Mem_reg[75][4]  ( .D(n24731), .E(n6406), .CP(clk), .QN(n27054) );
  EDFD1 \Mem_reg[74][4]  ( .D(n24731), .E(n6405), .CP(clk), .QN(n5718) );
  EDFD1 \Mem_reg[73][4]  ( .D(n24731), .E(n6404), .CP(clk), .QN(n27055) );
  EDFD1 \Mem_reg[72][4]  ( .D(n24731), .E(n6403), .CP(clk), .QN(n5622) );
  EDFD1 \Mem_reg[71][4]  ( .D(n24731), .E(n6402), .CP(clk), .QN(n5574) );
  EDFD1 \Mem_reg[70][4]  ( .D(n24731), .E(n6401), .CP(clk), .QN(n5526) );
  EDFD1 \Mem_reg[69][4]  ( .D(n24731), .E(n6400), .CP(clk), .QN(n5478) );
  EDFD1 \Mem_reg[68][4]  ( .D(n24731), .E(n6399), .CP(clk), .QN(n5430) );
  EDFD1 \Mem_reg[67][4]  ( .D(n24731), .E(n6398), .CP(clk), .QN(n5382) );
  EDFD1 \Mem_reg[66][4]  ( .D(n24731), .E(n6397), .CP(clk), .QN(n5334) );
  EDFD1 \Mem_reg[65][4]  ( .D(n24731), .E(n6396), .CP(clk), .QN(n15465) );
  EDFD1 \Mem_reg[64][4]  ( .D(n24731), .E(n6395), .CP(clk), .QN(n5238) );
  EDFD1 \Mem_reg[63][4]  ( .D(n24731), .E(n6456), .CP(clk), .QN(n5190) );
  EDFD1 \Mem_reg[62][4]  ( .D(n24731), .E(n6455), .CP(clk), .QN(n5142) );
  EDFD1 \Mem_reg[61][4]  ( .D(n24731), .E(n6454), .CP(clk), .QN(n17939) );
  EDFD1 \Mem_reg[60][4]  ( .D(n24731), .E(n6453), .CP(clk), .QN(n17938) );
  EDFD1 \Mem_reg[59][4]  ( .D(n24731), .E(n6452), .CP(clk), .QN(n4998) );
  EDFD1 \Mem_reg[58][4]  ( .D(n24731), .E(n6451), .CP(clk), .QN(n4950) );
  EDFD1 \Mem_reg[57][4]  ( .D(n24731), .E(n6450), .CP(clk), .QN(n4902) );
  EDFD1 \Mem_reg[56][4]  ( .D(n24731), .E(n6449), .CP(clk), .QN(n4854) );
  EDFD1 \Mem_reg[55][4]  ( .D(n24731), .E(n6448), .CP(clk), .QN(n4806) );
  EDFD1 \Mem_reg[54][4]  ( .D(n24731), .E(n6447), .CP(clk), .QN(n15464) );
  EDFD1 \Mem_reg[53][4]  ( .D(n24731), .E(n6446), .CP(clk), .QN(n4710) );
  EDFD1 \Mem_reg[52][4]  ( .D(n24731), .E(n6445), .CP(clk), .Q(n27052) );
  EDFD1 \Mem_reg[51][4]  ( .D(n24731), .E(n6444), .CP(clk), .QN(n4614) );
  EDFD1 \Mem_reg[50][4]  ( .D(n24731), .E(n6443), .CP(clk), .QN(n4566) );
  EDFD1 \Mem_reg[49][4]  ( .D(n24731), .E(n6442), .CP(clk), .QN(n4518) );
  EDFD1 \Mem_reg[48][4]  ( .D(n24731), .E(n6441), .CP(clk), .QN(n4470) );
  EDFD1 \Mem_reg[47][4]  ( .D(n24731), .E(n6440), .CP(clk), .QN(n4422) );
  EDFD1 \Mem_reg[46][4]  ( .D(n24731), .E(n6439), .CP(clk), .QN(n4374) );
  EDFD1 \Mem_reg[43][4]  ( .D(n24731), .E(n6438), .CP(clk), .QN(n4326) );
  EDFD1 \Mem_reg[42][4]  ( .D(n24731), .E(n6437), .CP(clk), .QN(n4278) );
  EDFD1 \Mem_reg[41][4]  ( .D(n24731), .E(n6436), .CP(clk), .QN(n4230) );
  EDFD1 \Mem_reg[40][4]  ( .D(n24731), .E(n6435), .CP(clk), .QN(n4182) );
  EDFD1 \Mem_reg[39][4]  ( .D(n24731), .E(n6434), .CP(clk), .QN(n4134) );
  EDFD1 \Mem_reg[38][4]  ( .D(n24731), .E(n6433), .CP(clk), .QN(n4086) );
  EDFD1 \Mem_reg[37][4]  ( .D(n24731), .E(n6432), .CP(clk), .QN(n4038) );
  EDFD1 \Mem_reg[36][4]  ( .D(n24731), .E(n6431), .CP(clk), .QN(n3990) );
  EDFD1 \Mem_reg[35][4]  ( .D(n24731), .E(n6430), .CP(clk), .QN(n3942) );
  EDFD1 \Mem_reg[34][4]  ( .D(n24731), .E(n6429), .CP(clk), .QN(n3894) );
  EDFD1 \Mem_reg[33][4]  ( .D(n24731), .E(n6428), .CP(clk), .QN(n3846) );
  EDFD1 \Mem_reg[32][4]  ( .D(n24731), .E(n6427), .CP(clk), .QN(n3798) );
  EDFD1 \Mem_reg[31][4]  ( .D(n24731), .E(n6426), .CP(clk), .QN(n3750) );
  EDFD1 \Mem_reg[30][4]  ( .D(n24731), .E(n6425), .CP(clk), .QN(n3702) );
  EDFD1 \Mem_reg[29][4]  ( .D(n24731), .E(n6424), .CP(clk), .QN(n3654) );
  EDFD1 \Mem_reg[28][4]  ( .D(n24731), .E(n6423), .CP(clk), .QN(n3606) );
  EDFD1 \Mem_reg[27][4]  ( .D(n24731), .E(n6422), .CP(clk), .QN(n3558) );
  EDFD1 \Mem_reg[26][4]  ( .D(n24731), .E(n6421), .CP(clk), .QN(n3510) );
  EDFD1 \Mem_reg[25][4]  ( .D(n24731), .E(n6420), .CP(clk), .QN(n3462) );
  EDFD1 \Mem_reg[24][4]  ( .D(n24731), .E(n6463), .CP(clk), .QN(n3414) );
  EDFD1 \Mem_reg[23][4]  ( .D(n24731), .E(n6464), .CP(clk), .QN(n3366) );
  EDFD1 \Mem_reg[22][4]  ( .D(n24731), .E(n6465), .CP(clk), .QN(n3318) );
  EDFD1 \Mem_reg[21][4]  ( .D(n24731), .E(n6466), .CP(clk), .QN(n3270) );
  EDFD1 \Mem_reg[20][4]  ( .D(n24731), .E(n6467), .CP(clk), .QN(n3222) );
  EDFD1 \Mem_reg[19][4]  ( .D(n24731), .E(n6468), .CP(clk), .QN(n3174) );
  EDFD1 \Mem_reg[18][4]  ( .D(n24731), .E(n6469), .CP(clk), .QN(n3126) );
  EDFD1 \Mem_reg[17][4]  ( .D(n24731), .E(n6470), .CP(clk), .QN(n3078) );
  EDFD1 \Mem_reg[16][4]  ( .D(n24731), .E(n6471), .CP(clk), .QN(n3030) );
  EDFD1 \Mem_reg[15][4]  ( .D(n24731), .E(n6472), .CP(clk), .QN(n2982) );
  EDFD1 \Mem_reg[14][4]  ( .D(n24731), .E(n24720), .CP(clk), .QN(n2934) );
  EDFD1 \Mem_reg[13][4]  ( .D(n24731), .E(n24709), .CP(clk), .QN(n2886) );
  EDFD1 \Mem_reg[12][4]  ( .D(n24731), .E(n24717), .CP(clk), .QN(n2838) );
  EDFD1 \Mem_reg[11][4]  ( .D(n24731), .E(n24707), .CP(clk), .QN(n2790) );
  EDFD1 \Mem_reg[10][4]  ( .D(n24731), .E(n6477), .CP(clk), .QN(n2742) );
  EDFD1 \Mem_reg[9][4]  ( .D(n24731), .E(n24708), .CP(clk), .QN(n2694) );
  EDFD1 \Mem_reg[8][4]  ( .D(n24731), .E(n15642), .CP(clk), .QN(n2646) );
  EDFD1 \Mem_reg[7][4]  ( .D(n24731), .E(n24718), .CP(clk), .QN(n2598) );
  EDFD1 \Mem_reg[6][4]  ( .D(n24731), .E(n24716), .CP(clk), .QN(n2550) );
  EDFD1 \Mem_reg[5][4]  ( .D(n24731), .E(n24719), .CP(clk), .QN(n2502) );
  EDFD1 \Mem_reg[4][4]  ( .D(n24731), .E(n24706), .CP(clk), .QN(n2454) );
  EDFD1 \Mem_reg[3][4]  ( .D(n24731), .E(n24721), .CP(clk), .QN(n2406) );
  EDFD1 \Mem_reg[2][4]  ( .D(n24731), .E(n6460), .CP(clk), .QN(n2358) );
  EDFD1 \Mem_reg[1][4]  ( .D(n24731), .E(n24703), .CP(clk), .QN(n2310) );
  EDFD1 \Mem_reg[0][4]  ( .D(n24731), .E(n24705), .CP(clk), .QN(n2262) );
  EDFD1 \Mem_reg[88][3]  ( .D(n24729), .E(n6419), .CP(clk), .Q(n27049) );
  EDFD1 \Mem_reg[87][3]  ( .D(n24729), .E(n6418), .CP(clk), .QN(n6343) );
  EDFD1 \Mem_reg[86][3]  ( .D(n24729), .E(n6417), .CP(clk), .QN(n24568) );
  EDFD1 \Mem_reg[85][3]  ( .D(n24729), .E(n6416), .CP(clk), .QN(n6247) );
  EDFD1 \Mem_reg[84][3]  ( .D(n24729), .E(n6415), .CP(clk), .QN(n6199) );
  EDFD1 \Mem_reg[83][3]  ( .D(n24729), .E(n6414), .CP(clk), .QN(n6151) );
  EDFD1 \Mem_reg[82][3]  ( .D(n24729), .E(n6413), .CP(clk), .QN(n6103) );
  EDFD1 \Mem_reg[81][3]  ( .D(n24729), .E(n6412), .CP(clk), .QN(n6055) );
  EDFD1 \Mem_reg[80][3]  ( .D(n24729), .E(n6411), .CP(clk), .QN(n6007) );
  EDFD1 \Mem_reg[79][3]  ( .D(n24729), .E(n6410), .CP(clk), .QN(n5959) );
  EDFD1 \Mem_reg[78][3]  ( .D(n24729), .E(n6409), .CP(clk), .QN(n5911) );
  EDFD1 \Mem_reg[77][3]  ( .D(n24729), .E(n6408), .CP(clk), .QN(n5863) );
  EDFD1 \Mem_reg[76][3]  ( .D(n24729), .E(n6407), .CP(clk), .QN(n5815) );
  EDFD1 \Mem_reg[75][3]  ( .D(n24729), .E(n6406), .CP(clk), .QN(n27050) );
  EDFD1 \Mem_reg[74][3]  ( .D(n24729), .E(n6405), .CP(clk), .QN(n5719) );
  EDFD1 \Mem_reg[73][3]  ( .D(n24729), .E(n6404), .CP(clk), .QN(n27051) );
  EDFD1 \Mem_reg[72][3]  ( .D(n24729), .E(n6403), .CP(clk), .QN(n5623) );
  EDFD1 \Mem_reg[71][3]  ( .D(n24729), .E(n6402), .CP(clk), .QN(n5575) );
  EDFD1 \Mem_reg[70][3]  ( .D(n24729), .E(n6401), .CP(clk), .QN(n5527) );
  EDFD1 \Mem_reg[69][3]  ( .D(n24729), .E(n6400), .CP(clk), .QN(n5479) );
  EDFD1 \Mem_reg[68][3]  ( .D(n24729), .E(n6399), .CP(clk), .QN(n5431) );
  EDFD1 \Mem_reg[67][3]  ( .D(n24729), .E(n6398), .CP(clk), .QN(n5383) );
  EDFD1 \Mem_reg[66][3]  ( .D(n24729), .E(n6397), .CP(clk), .QN(n5335) );
  EDFD1 \Mem_reg[65][3]  ( .D(n24729), .E(n6396), .CP(clk), .QN(n15461) );
  EDFD1 \Mem_reg[64][3]  ( .D(n24729), .E(n6395), .CP(clk), .QN(n5239) );
  EDFD1 \Mem_reg[63][3]  ( .D(n24729), .E(n6456), .CP(clk), .QN(n5191) );
  EDFD1 \Mem_reg[62][3]  ( .D(n24729), .E(n6455), .CP(clk), .QN(n5143) );
  EDFD1 \Mem_reg[61][3]  ( .D(n24729), .E(n6454), .CP(clk), .QN(n17936) );
  EDFD1 \Mem_reg[60][3]  ( .D(n24729), .E(n6453), .CP(clk), .QN(n17935) );
  EDFD1 \Mem_reg[59][3]  ( .D(n24729), .E(n6452), .CP(clk), .QN(n4999) );
  EDFD1 \Mem_reg[58][3]  ( .D(n24729), .E(n6451), .CP(clk), .QN(n4951) );
  EDFD1 \Mem_reg[57][3]  ( .D(n24729), .E(n6450), .CP(clk), .QN(n4903) );
  EDFD1 \Mem_reg[56][3]  ( .D(n24729), .E(n6449), .CP(clk), .QN(n4855) );
  EDFD1 \Mem_reg[55][3]  ( .D(n24729), .E(n6448), .CP(clk), .QN(n4807) );
  EDFD1 \Mem_reg[54][3]  ( .D(n24729), .E(n6447), .CP(clk), .QN(n15460) );
  EDFD1 \Mem_reg[53][3]  ( .D(n24729), .E(n6446), .CP(clk), .QN(n4711) );
  EDFD1 \Mem_reg[52][3]  ( .D(n24729), .E(n6445), .CP(clk), .Q(n27048) );
  EDFD1 \Mem_reg[51][3]  ( .D(n24729), .E(n6444), .CP(clk), .QN(n4615) );
  EDFD1 \Mem_reg[50][3]  ( .D(n24729), .E(n6443), .CP(clk), .QN(n4567) );
  EDFD1 \Mem_reg[49][3]  ( .D(n24729), .E(n6442), .CP(clk), .QN(n4519) );
  EDFD1 \Mem_reg[48][3]  ( .D(n24729), .E(n6441), .CP(clk), .QN(n4471) );
  EDFD1 \Mem_reg[47][3]  ( .D(n24729), .E(n6440), .CP(clk), .QN(n4423) );
  EDFD1 \Mem_reg[46][3]  ( .D(n24729), .E(n6439), .CP(clk), .QN(n4375) );
  EDFD1 \Mem_reg[43][3]  ( .D(n24729), .E(n6438), .CP(clk), .QN(n4327) );
  EDFD1 \Mem_reg[42][3]  ( .D(n24729), .E(n6437), .CP(clk), .QN(n4279) );
  EDFD1 \Mem_reg[41][3]  ( .D(n24729), .E(n6436), .CP(clk), .QN(n4231) );
  EDFD1 \Mem_reg[40][3]  ( .D(n24729), .E(n6435), .CP(clk), .QN(n4183) );
  EDFD1 \Mem_reg[39][3]  ( .D(n24729), .E(n6434), .CP(clk), .QN(n4135) );
  EDFD1 \Mem_reg[38][3]  ( .D(n24729), .E(n6433), .CP(clk), .QN(n4087) );
  EDFD1 \Mem_reg[37][3]  ( .D(n24729), .E(n6432), .CP(clk), .QN(n4039) );
  EDFD1 \Mem_reg[36][3]  ( .D(n24729), .E(n6431), .CP(clk), .QN(n3991) );
  EDFD1 \Mem_reg[35][3]  ( .D(n24729), .E(n6430), .CP(clk), .QN(n3943) );
  EDFD1 \Mem_reg[34][3]  ( .D(n24729), .E(n6429), .CP(clk), .QN(n3895) );
  EDFD1 \Mem_reg[33][3]  ( .D(n24729), .E(n6428), .CP(clk), .QN(n3847) );
  EDFD1 \Mem_reg[32][3]  ( .D(n24729), .E(n6427), .CP(clk), .QN(n3799) );
  EDFD1 \Mem_reg[31][3]  ( .D(n24729), .E(n6426), .CP(clk), .QN(n3751) );
  EDFD1 \Mem_reg[30][3]  ( .D(n24729), .E(n6425), .CP(clk), .QN(n3703) );
  EDFD1 \Mem_reg[29][3]  ( .D(n24729), .E(n6424), .CP(clk), .QN(n3655) );
  EDFD1 \Mem_reg[28][3]  ( .D(n24729), .E(n6423), .CP(clk), .QN(n3607) );
  EDFD1 \Mem_reg[27][3]  ( .D(n24729), .E(n6422), .CP(clk), .QN(n3559) );
  EDFD1 \Mem_reg[26][3]  ( .D(n24729), .E(n6421), .CP(clk), .QN(n3511) );
  EDFD1 \Mem_reg[25][3]  ( .D(n24729), .E(n6420), .CP(clk), .QN(n3463) );
  EDFD1 \Mem_reg[24][3]  ( .D(n24729), .E(n6463), .CP(clk), .QN(n3415) );
  EDFD1 \Mem_reg[23][3]  ( .D(n24729), .E(n6464), .CP(clk), .QN(n3367) );
  EDFD1 \Mem_reg[22][3]  ( .D(n24729), .E(n6465), .CP(clk), .QN(n3319) );
  EDFD1 \Mem_reg[21][3]  ( .D(n24729), .E(n6466), .CP(clk), .QN(n3271) );
  EDFD1 \Mem_reg[20][3]  ( .D(n24729), .E(n6467), .CP(clk), .QN(n3223) );
  EDFD1 \Mem_reg[19][3]  ( .D(n24729), .E(n6468), .CP(clk), .QN(n3175) );
  EDFD1 \Mem_reg[18][3]  ( .D(n24729), .E(n6469), .CP(clk), .QN(n3127) );
  EDFD1 \Mem_reg[17][3]  ( .D(n24729), .E(n6470), .CP(clk), .QN(n3079) );
  EDFD1 \Mem_reg[16][3]  ( .D(n24729), .E(n6471), .CP(clk), .QN(n3031) );
  EDFD1 \Mem_reg[15][3]  ( .D(n24729), .E(n6472), .CP(clk), .QN(n2983) );
  EDFD1 \Mem_reg[14][3]  ( .D(n24729), .E(n24720), .CP(clk), .QN(n2935) );
  EDFD1 \Mem_reg[13][3]  ( .D(n24729), .E(n24709), .CP(clk), .QN(n2887) );
  EDFD1 \Mem_reg[12][3]  ( .D(n24729), .E(n24717), .CP(clk), .QN(n2839) );
  EDFD1 \Mem_reg[11][3]  ( .D(n24729), .E(n24707), .CP(clk), .QN(n2791) );
  EDFD1 \Mem_reg[10][3]  ( .D(n24729), .E(n6477), .CP(clk), .QN(n2743) );
  EDFD1 \Mem_reg[9][3]  ( .D(n24729), .E(n24708), .CP(clk), .QN(n2695) );
  EDFD1 \Mem_reg[8][3]  ( .D(n24729), .E(n15642), .CP(clk), .QN(n2647) );
  EDFD1 \Mem_reg[7][3]  ( .D(n24729), .E(n24718), .CP(clk), .QN(n2599) );
  EDFD1 \Mem_reg[6][3]  ( .D(n24729), .E(n24716), .CP(clk), .QN(n2551) );
  EDFD1 \Mem_reg[5][3]  ( .D(n24729), .E(n24719), .CP(clk), .QN(n2503) );
  EDFD1 \Mem_reg[4][3]  ( .D(n24729), .E(n24706), .CP(clk), .QN(n2455) );
  EDFD1 \Mem_reg[3][3]  ( .D(n24729), .E(n24721), .CP(clk), .QN(n2407) );
  EDFD1 \Mem_reg[2][3]  ( .D(n24729), .E(n6460), .CP(clk), .QN(n2359) );
  EDFD1 \Mem_reg[1][3]  ( .D(n24729), .E(n24703), .CP(clk), .QN(n2311) );
  EDFD1 \Mem_reg[0][3]  ( .D(n24729), .E(n24705), .CP(clk), .QN(n2263) );
  EDFD1 \Mem_reg[88][2]  ( .D(n24727), .E(n6419), .CP(clk), .Q(n27045) );
  EDFD1 \Mem_reg[87][2]  ( .D(n24727), .E(n6418), .CP(clk), .QN(n6344) );
  EDFD1 \Mem_reg[86][2]  ( .D(n24727), .E(n6417), .CP(clk), .QN(n24565) );
  EDFD1 \Mem_reg[85][2]  ( .D(n24727), .E(n6416), .CP(clk), .QN(n6248) );
  EDFD1 \Mem_reg[84][2]  ( .D(n24727), .E(n6415), .CP(clk), .QN(n6200) );
  EDFD1 \Mem_reg[83][2]  ( .D(n24727), .E(n6414), .CP(clk), .QN(n6152) );
  EDFD1 \Mem_reg[82][2]  ( .D(n24727), .E(n6413), .CP(clk), .QN(n6104) );
  EDFD1 \Mem_reg[81][2]  ( .D(n24727), .E(n6412), .CP(clk), .QN(n6056) );
  EDFD1 \Mem_reg[80][2]  ( .D(n24727), .E(n6411), .CP(clk), .QN(n6008) );
  EDFD1 \Mem_reg[79][2]  ( .D(n24727), .E(n6410), .CP(clk), .QN(n5960) );
  EDFD1 \Mem_reg[78][2]  ( .D(n24727), .E(n6409), .CP(clk), .QN(n5912) );
  EDFD1 \Mem_reg[77][2]  ( .D(n24727), .E(n6408), .CP(clk), .QN(n5864) );
  EDFD1 \Mem_reg[76][2]  ( .D(n24727), .E(n6407), .CP(clk), .QN(n5816) );
  EDFD1 \Mem_reg[75][2]  ( .D(n24727), .E(n6406), .CP(clk), .QN(n27046) );
  EDFD1 \Mem_reg[74][2]  ( .D(n24727), .E(n6405), .CP(clk), .QN(n5720) );
  EDFD1 \Mem_reg[73][2]  ( .D(n24727), .E(n6404), .CP(clk), .QN(n27047) );
  EDFD1 \Mem_reg[72][2]  ( .D(n24727), .E(n6403), .CP(clk), .QN(n5624) );
  EDFD1 \Mem_reg[71][2]  ( .D(n24727), .E(n6402), .CP(clk), .QN(n5576) );
  EDFD1 \Mem_reg[70][2]  ( .D(n24727), .E(n6401), .CP(clk), .QN(n5528) );
  EDFD1 \Mem_reg[69][2]  ( .D(n24727), .E(n6400), .CP(clk), .QN(n5480) );
  EDFD1 \Mem_reg[68][2]  ( .D(n24727), .E(n6399), .CP(clk), .QN(n5432) );
  EDFD1 \Mem_reg[67][2]  ( .D(n24727), .E(n6398), .CP(clk), .QN(n5384) );
  EDFD1 \Mem_reg[66][2]  ( .D(n24727), .E(n6397), .CP(clk), .QN(n5336) );
  EDFD1 \Mem_reg[65][2]  ( .D(n24727), .E(n6396), .CP(clk), .QN(n15457) );
  EDFD1 \Mem_reg[64][2]  ( .D(n24727), .E(n6395), .CP(clk), .QN(n5240) );
  EDFD1 \Mem_reg[63][2]  ( .D(n24727), .E(n6456), .CP(clk), .QN(n5192) );
  EDFD1 \Mem_reg[62][2]  ( .D(n24727), .E(n6455), .CP(clk), .QN(n5144) );
  EDFD1 \Mem_reg[61][2]  ( .D(n24727), .E(n6454), .CP(clk), .QN(n17933) );
  EDFD1 \Mem_reg[60][2]  ( .D(n24727), .E(n6453), .CP(clk), .QN(n17932) );
  EDFD1 \Mem_reg[59][2]  ( .D(n24727), .E(n6452), .CP(clk), .QN(n5000) );
  EDFD1 \Mem_reg[58][2]  ( .D(n24727), .E(n6451), .CP(clk), .QN(n4952) );
  EDFD1 \Mem_reg[57][2]  ( .D(n24727), .E(n6450), .CP(clk), .QN(n4904) );
  EDFD1 \Mem_reg[56][2]  ( .D(n24727), .E(n6449), .CP(clk), .QN(n4856) );
  EDFD1 \Mem_reg[55][2]  ( .D(n24727), .E(n6448), .CP(clk), .QN(n4808) );
  EDFD1 \Mem_reg[54][2]  ( .D(n24727), .E(n6447), .CP(clk), .QN(n15456) );
  EDFD1 \Mem_reg[53][2]  ( .D(n24727), .E(n6446), .CP(clk), .QN(n4712) );
  EDFD1 \Mem_reg[52][2]  ( .D(n24727), .E(n6445), .CP(clk), .Q(n27044) );
  EDFD1 \Mem_reg[51][2]  ( .D(n24727), .E(n6444), .CP(clk), .QN(n4616) );
  EDFD1 \Mem_reg[50][2]  ( .D(n24727), .E(n6443), .CP(clk), .QN(n4568) );
  EDFD1 \Mem_reg[49][2]  ( .D(n24727), .E(n6442), .CP(clk), .QN(n4520) );
  EDFD1 \Mem_reg[48][2]  ( .D(n24727), .E(n6441), .CP(clk), .QN(n4472) );
  EDFD1 \Mem_reg[47][2]  ( .D(n24727), .E(n6440), .CP(clk), .QN(n4424) );
  EDFD1 \Mem_reg[46][2]  ( .D(n24727), .E(n6439), .CP(clk), .QN(n4376) );
  EDFD1 \Mem_reg[43][2]  ( .D(n24727), .E(n6438), .CP(clk), .QN(n4328) );
  EDFD1 \Mem_reg[42][2]  ( .D(n24727), .E(n6437), .CP(clk), .QN(n4280) );
  EDFD1 \Mem_reg[41][2]  ( .D(n24727), .E(n6436), .CP(clk), .QN(n4232) );
  EDFD1 \Mem_reg[40][2]  ( .D(n24727), .E(n6435), .CP(clk), .QN(n4184) );
  EDFD1 \Mem_reg[39][2]  ( .D(n24727), .E(n6434), .CP(clk), .QN(n4136) );
  EDFD1 \Mem_reg[38][2]  ( .D(n24727), .E(n6433), .CP(clk), .QN(n4088) );
  EDFD1 \Mem_reg[37][2]  ( .D(n24727), .E(n6432), .CP(clk), .QN(n4040) );
  EDFD1 \Mem_reg[36][2]  ( .D(n24727), .E(n6431), .CP(clk), .QN(n3992) );
  EDFD1 \Mem_reg[35][2]  ( .D(n24727), .E(n6430), .CP(clk), .QN(n3944) );
  EDFD1 \Mem_reg[34][2]  ( .D(n24727), .E(n6429), .CP(clk), .QN(n3896) );
  EDFD1 \Mem_reg[33][2]  ( .D(n24727), .E(n6428), .CP(clk), .QN(n3848) );
  EDFD1 \Mem_reg[32][2]  ( .D(n24727), .E(n6427), .CP(clk), .QN(n3800) );
  EDFD1 \Mem_reg[31][2]  ( .D(n24727), .E(n6426), .CP(clk), .QN(n3752) );
  EDFD1 \Mem_reg[30][2]  ( .D(n24727), .E(n6425), .CP(clk), .QN(n3704) );
  EDFD1 \Mem_reg[29][2]  ( .D(n24727), .E(n6424), .CP(clk), .QN(n3656) );
  EDFD1 \Mem_reg[28][2]  ( .D(n24727), .E(n6423), .CP(clk), .QN(n3608) );
  EDFD1 \Mem_reg[27][2]  ( .D(n24727), .E(n6422), .CP(clk), .QN(n3560) );
  EDFD1 \Mem_reg[26][2]  ( .D(n24727), .E(n6421), .CP(clk), .QN(n3512) );
  EDFD1 \Mem_reg[25][2]  ( .D(n24727), .E(n6420), .CP(clk), .QN(n3464) );
  EDFD1 \Mem_reg[24][2]  ( .D(n24727), .E(n6463), .CP(clk), .QN(n3416) );
  EDFD1 \Mem_reg[23][2]  ( .D(n24727), .E(n6464), .CP(clk), .QN(n3368) );
  EDFD1 \Mem_reg[22][2]  ( .D(n24727), .E(n6465), .CP(clk), .QN(n3320) );
  EDFD1 \Mem_reg[21][2]  ( .D(n24727), .E(n6466), .CP(clk), .QN(n3272) );
  EDFD1 \Mem_reg[20][2]  ( .D(n24727), .E(n6467), .CP(clk), .QN(n3224) );
  EDFD1 \Mem_reg[19][2]  ( .D(n24727), .E(n6468), .CP(clk), .QN(n3176) );
  EDFD1 \Mem_reg[18][2]  ( .D(n24727), .E(n6469), .CP(clk), .QN(n3128) );
  EDFD1 \Mem_reg[17][2]  ( .D(n24727), .E(n6470), .CP(clk), .QN(n3080) );
  EDFD1 \Mem_reg[16][2]  ( .D(n24727), .E(n6471), .CP(clk), .QN(n3032) );
  EDFD1 \Mem_reg[15][2]  ( .D(n24727), .E(n6472), .CP(clk), .QN(n2984) );
  EDFD1 \Mem_reg[14][2]  ( .D(n24727), .E(n24720), .CP(clk), .QN(n2936) );
  EDFD1 \Mem_reg[13][2]  ( .D(n24727), .E(n24709), .CP(clk), .QN(n2888) );
  EDFD1 \Mem_reg[12][2]  ( .D(n24727), .E(n24717), .CP(clk), .QN(n2840) );
  EDFD1 \Mem_reg[11][2]  ( .D(n24727), .E(n24707), .CP(clk), .QN(n2792) );
  EDFD1 \Mem_reg[10][2]  ( .D(n24727), .E(n6477), .CP(clk), .QN(n2744) );
  EDFD1 \Mem_reg[9][2]  ( .D(n24727), .E(n24708), .CP(clk), .QN(n2696) );
  EDFD1 \Mem_reg[8][2]  ( .D(n24727), .E(n15642), .CP(clk), .QN(n2648) );
  EDFD1 \Mem_reg[7][2]  ( .D(n24727), .E(n24718), .CP(clk), .QN(n2600) );
  EDFD1 \Mem_reg[6][2]  ( .D(n24727), .E(n24716), .CP(clk), .QN(n2552) );
  EDFD1 \Mem_reg[5][2]  ( .D(n24727), .E(n24719), .CP(clk), .QN(n2504) );
  EDFD1 \Mem_reg[4][2]  ( .D(n24727), .E(n24706), .CP(clk), .QN(n2456) );
  EDFD1 \Mem_reg[3][2]  ( .D(n24727), .E(n24721), .CP(clk), .QN(n2408) );
  EDFD1 \Mem_reg[2][2]  ( .D(n24727), .E(n6460), .CP(clk), .QN(n2360) );
  EDFD1 \Mem_reg[1][2]  ( .D(n24727), .E(n24703), .CP(clk), .QN(n2312) );
  EDFD1 \Mem_reg[0][2]  ( .D(n24727), .E(n24705), .CP(clk), .QN(n2264) );
  EDFD1 \Mem_reg[88][1]  ( .D(n24725), .E(n6419), .CP(clk), .Q(n27041) );
  EDFD1 \Mem_reg[87][1]  ( .D(n24725), .E(n6418), .CP(clk), .QN(n6345) );
  EDFD1 \Mem_reg[86][1]  ( .D(n24725), .E(n6417), .CP(clk), .QN(n24562) );
  EDFD1 \Mem_reg[85][1]  ( .D(n24725), .E(n6416), .CP(clk), .QN(n6249) );
  EDFD1 \Mem_reg[84][1]  ( .D(n24725), .E(n6415), .CP(clk), .QN(n6201) );
  EDFD1 \Mem_reg[83][1]  ( .D(n24725), .E(n6414), .CP(clk), .QN(n6153) );
  EDFD1 \Mem_reg[82][1]  ( .D(n24725), .E(n6413), .CP(clk), .QN(n6105) );
  EDFD1 \Mem_reg[81][1]  ( .D(n24725), .E(n6412), .CP(clk), .QN(n6057) );
  EDFD1 \Mem_reg[80][1]  ( .D(n24725), .E(n6411), .CP(clk), .QN(n6009) );
  EDFD1 \Mem_reg[79][1]  ( .D(n24725), .E(n6410), .CP(clk), .QN(n5961) );
  EDFD1 \Mem_reg[78][1]  ( .D(n24725), .E(n6409), .CP(clk), .QN(n5913) );
  EDFD1 \Mem_reg[77][1]  ( .D(n24725), .E(n6408), .CP(clk), .QN(n5865) );
  EDFD1 \Mem_reg[76][1]  ( .D(n24725), .E(n6407), .CP(clk), .QN(n5817) );
  EDFD1 \Mem_reg[75][1]  ( .D(n24725), .E(n6406), .CP(clk), .QN(n27042) );
  EDFD1 \Mem_reg[74][1]  ( .D(n24725), .E(n6405), .CP(clk), .QN(n5721) );
  EDFD1 \Mem_reg[73][1]  ( .D(n24725), .E(n6404), .CP(clk), .QN(n27043) );
  EDFD1 \Mem_reg[72][1]  ( .D(n24725), .E(n6403), .CP(clk), .QN(n5625) );
  EDFD1 \Mem_reg[71][1]  ( .D(n24725), .E(n6402), .CP(clk), .QN(n5577) );
  EDFD1 \Mem_reg[70][1]  ( .D(n24725), .E(n6401), .CP(clk), .QN(n5529) );
  EDFD1 \Mem_reg[69][1]  ( .D(n24725), .E(n6400), .CP(clk), .QN(n5481) );
  EDFD1 \Mem_reg[68][1]  ( .D(n24725), .E(n6399), .CP(clk), .QN(n5433) );
  EDFD1 \Mem_reg[67][1]  ( .D(n24725), .E(n6398), .CP(clk), .QN(n5385) );
  EDFD1 \Mem_reg[66][1]  ( .D(n24725), .E(n6397), .CP(clk), .QN(n5337) );
  EDFD1 \Mem_reg[65][1]  ( .D(n24725), .E(n6396), .CP(clk), .QN(n15453) );
  EDFD1 \Mem_reg[64][1]  ( .D(n24725), .E(n6395), .CP(clk), .QN(n5241) );
  EDFD1 \Mem_reg[63][1]  ( .D(n24725), .E(n6456), .CP(clk), .QN(n5193) );
  EDFD1 \Mem_reg[62][1]  ( .D(n24725), .E(n6455), .CP(clk), .QN(n5145) );
  EDFD1 \Mem_reg[61][1]  ( .D(n24725), .E(n6454), .CP(clk), .QN(n17930) );
  EDFD1 \Mem_reg[60][1]  ( .D(n24725), .E(n6453), .CP(clk), .QN(n17929) );
  EDFD1 \Mem_reg[59][1]  ( .D(n24725), .E(n6452), .CP(clk), .QN(n5001) );
  EDFD1 \Mem_reg[58][1]  ( .D(n24725), .E(n6451), .CP(clk), .QN(n4953) );
  EDFD1 \Mem_reg[57][1]  ( .D(n24725), .E(n6450), .CP(clk), .QN(n4905) );
  EDFD1 \Mem_reg[56][1]  ( .D(n24725), .E(n6449), .CP(clk), .QN(n4857) );
  EDFD1 \Mem_reg[55][1]  ( .D(n24725), .E(n6448), .CP(clk), .QN(n4809) );
  EDFD1 \Mem_reg[54][1]  ( .D(n24725), .E(n6447), .CP(clk), .QN(n15452) );
  EDFD1 \Mem_reg[53][1]  ( .D(n24725), .E(n6446), .CP(clk), .QN(n4713) );
  EDFD1 \Mem_reg[52][1]  ( .D(n24725), .E(n6445), .CP(clk), .Q(n27040) );
  EDFD1 \Mem_reg[51][1]  ( .D(n24725), .E(n6444), .CP(clk), .QN(n4617) );
  EDFD1 \Mem_reg[50][1]  ( .D(n24725), .E(n6443), .CP(clk), .QN(n4569) );
  EDFD1 \Mem_reg[49][1]  ( .D(n24725), .E(n6442), .CP(clk), .QN(n4521) );
  EDFD1 \Mem_reg[48][1]  ( .D(n24725), .E(n6441), .CP(clk), .QN(n4473) );
  EDFD1 \Mem_reg[47][1]  ( .D(n24725), .E(n6440), .CP(clk), .QN(n4425) );
  EDFD1 \Mem_reg[46][1]  ( .D(n24725), .E(n6439), .CP(clk), .QN(n4377) );
  EDFD1 \Mem_reg[43][1]  ( .D(n24725), .E(n6438), .CP(clk), .QN(n4329) );
  EDFD1 \Mem_reg[42][1]  ( .D(n24725), .E(n6437), .CP(clk), .QN(n4281) );
  EDFD1 \Mem_reg[41][1]  ( .D(n24725), .E(n6436), .CP(clk), .QN(n4233) );
  EDFD1 \Mem_reg[40][1]  ( .D(n24725), .E(n6435), .CP(clk), .QN(n4185) );
  EDFD1 \Mem_reg[39][1]  ( .D(n24725), .E(n6434), .CP(clk), .QN(n4137) );
  EDFD1 \Mem_reg[38][1]  ( .D(n24725), .E(n6433), .CP(clk), .QN(n4089) );
  EDFD1 \Mem_reg[37][1]  ( .D(n24725), .E(n6432), .CP(clk), .QN(n4041) );
  EDFD1 \Mem_reg[36][1]  ( .D(n24725), .E(n6431), .CP(clk), .QN(n3993) );
  EDFD1 \Mem_reg[35][1]  ( .D(n24725), .E(n6430), .CP(clk), .QN(n3945) );
  EDFD1 \Mem_reg[34][1]  ( .D(n24725), .E(n6429), .CP(clk), .QN(n3897) );
  EDFD1 \Mem_reg[33][1]  ( .D(n24725), .E(n6428), .CP(clk), .QN(n3849) );
  EDFD1 \Mem_reg[32][1]  ( .D(n24725), .E(n6427), .CP(clk), .QN(n3801) );
  EDFD1 \Mem_reg[31][1]  ( .D(n24725), .E(n6426), .CP(clk), .QN(n3753) );
  EDFD1 \Mem_reg[30][1]  ( .D(n24725), .E(n6425), .CP(clk), .QN(n3705) );
  EDFD1 \Mem_reg[29][1]  ( .D(n24725), .E(n6424), .CP(clk), .QN(n3657) );
  EDFD1 \Mem_reg[28][1]  ( .D(n24725), .E(n6423), .CP(clk), .QN(n3609) );
  EDFD1 \Mem_reg[27][1]  ( .D(n24725), .E(n6422), .CP(clk), .QN(n3561) );
  EDFD1 \Mem_reg[26][1]  ( .D(n24725), .E(n6421), .CP(clk), .QN(n3513) );
  EDFD1 \Mem_reg[25][1]  ( .D(n24725), .E(n6420), .CP(clk), .QN(n3465) );
  EDFD1 \Mem_reg[24][1]  ( .D(n24725), .E(n6463), .CP(clk), .QN(n3417) );
  EDFD1 \Mem_reg[23][1]  ( .D(n24725), .E(n6464), .CP(clk), .QN(n3369) );
  EDFD1 \Mem_reg[22][1]  ( .D(n24725), .E(n6465), .CP(clk), .QN(n3321) );
  EDFD1 \Mem_reg[21][1]  ( .D(n24725), .E(n6466), .CP(clk), .QN(n3273) );
  EDFD1 \Mem_reg[20][1]  ( .D(n24725), .E(n6467), .CP(clk), .QN(n3225) );
  EDFD1 \Mem_reg[19][1]  ( .D(n24725), .E(n6468), .CP(clk), .QN(n3177) );
  EDFD1 \Mem_reg[18][1]  ( .D(n24725), .E(n6469), .CP(clk), .QN(n3129) );
  EDFD1 \Mem_reg[17][1]  ( .D(n24725), .E(n6470), .CP(clk), .QN(n3081) );
  EDFD1 \Mem_reg[16][1]  ( .D(n24725), .E(n6471), .CP(clk), .QN(n3033) );
  EDFD1 \Mem_reg[15][1]  ( .D(n24725), .E(n6472), .CP(clk), .QN(n2985) );
  EDFD1 \Mem_reg[14][1]  ( .D(n24725), .E(n24720), .CP(clk), .QN(n2937) );
  EDFD1 \Mem_reg[13][1]  ( .D(n24725), .E(n24709), .CP(clk), .QN(n2889) );
  EDFD1 \Mem_reg[12][1]  ( .D(n24725), .E(n24717), .CP(clk), .QN(n2841) );
  EDFD1 \Mem_reg[11][1]  ( .D(n24725), .E(n24707), .CP(clk), .QN(n2793) );
  EDFD1 \Mem_reg[10][1]  ( .D(n24725), .E(n6477), .CP(clk), .QN(n2745) );
  EDFD1 \Mem_reg[9][1]  ( .D(n24725), .E(n24708), .CP(clk), .QN(n2697) );
  EDFD1 \Mem_reg[8][1]  ( .D(n24725), .E(n15642), .CP(clk), .QN(n2649) );
  EDFD1 \Mem_reg[7][1]  ( .D(n24725), .E(n24718), .CP(clk), .QN(n2601) );
  EDFD1 \Mem_reg[6][1]  ( .D(n24725), .E(n24716), .CP(clk), .QN(n2553) );
  EDFD1 \Mem_reg[5][1]  ( .D(n24725), .E(n24719), .CP(clk), .QN(n2505) );
  EDFD1 \Mem_reg[4][1]  ( .D(n24725), .E(n24706), .CP(clk), .QN(n2457) );
  EDFD1 \Mem_reg[3][1]  ( .D(n24725), .E(n24721), .CP(clk), .QN(n2409) );
  EDFD1 \Mem_reg[2][1]  ( .D(n24725), .E(n6460), .CP(clk), .QN(n2361) );
  EDFD1 \Mem_reg[1][1]  ( .D(n24725), .E(n24703), .CP(clk), .QN(n2313) );
  EDFD1 \Mem_reg[0][1]  ( .D(n24725), .E(n24705), .CP(clk), .QN(n2265) );
  EDFD1 \Mem_reg[88][0]  ( .D(n24723), .E(n6419), .CP(clk), .Q(n27037) );
  EDFD1 \Mem_reg[87][0]  ( .D(n24723), .E(n6418), .CP(clk), .QN(n6346) );
  EDFD1 \Mem_reg[86][0]  ( .D(n24723), .E(n6417), .CP(clk), .QN(n24559) );
  EDFD1 \Mem_reg[85][0]  ( .D(n24723), .E(n6416), .CP(clk), .QN(n6250) );
  EDFD1 \Mem_reg[84][0]  ( .D(n24723), .E(n6415), .CP(clk), .QN(n6202) );
  EDFD1 \Mem_reg[83][0]  ( .D(n24723), .E(n6414), .CP(clk), .QN(n6154) );
  EDFD1 \Mem_reg[82][0]  ( .D(n24723), .E(n6413), .CP(clk), .QN(n6106) );
  EDFD1 \Mem_reg[81][0]  ( .D(n24723), .E(n6412), .CP(clk), .QN(n6058) );
  EDFD1 \Mem_reg[80][0]  ( .D(n24723), .E(n6411), .CP(clk), .QN(n6010) );
  EDFD1 \Mem_reg[79][0]  ( .D(n24723), .E(n6410), .CP(clk), .QN(n5962) );
  EDFD1 \Mem_reg[78][0]  ( .D(n24723), .E(n6409), .CP(clk), .QN(n5914) );
  EDFD1 \Mem_reg[77][0]  ( .D(n24723), .E(n6408), .CP(clk), .QN(n5866) );
  EDFD1 \Mem_reg[76][0]  ( .D(n24723), .E(n6407), .CP(clk), .QN(n5818) );
  EDFD1 \Mem_reg[75][0]  ( .D(n24723), .E(n6406), .CP(clk), .QN(n27038) );
  EDFD1 \Mem_reg[74][0]  ( .D(n24723), .E(n6405), .CP(clk), .QN(n5722) );
  EDFD1 \Mem_reg[73][0]  ( .D(n24723), .E(n6404), .CP(clk), .QN(n27039) );
  EDFD1 \Mem_reg[72][0]  ( .D(n24723), .E(n6403), .CP(clk), .QN(n5626) );
  EDFD1 \Mem_reg[71][0]  ( .D(n24723), .E(n6402), .CP(clk), .QN(n5578) );
  EDFD1 \Mem_reg[70][0]  ( .D(n24723), .E(n6401), .CP(clk), .QN(n5530) );
  EDFD1 \Mem_reg[69][0]  ( .D(n24723), .E(n6400), .CP(clk), .QN(n5482) );
  EDFD1 \Mem_reg[68][0]  ( .D(n24723), .E(n6399), .CP(clk), .QN(n5434) );
  EDFD1 \Mem_reg[67][0]  ( .D(n24723), .E(n6398), .CP(clk), .QN(n5386) );
  EDFD1 \Mem_reg[66][0]  ( .D(n24723), .E(n6397), .CP(clk), .QN(n5338) );
  EDFD1 \Mem_reg[65][0]  ( .D(n24723), .E(n6396), .CP(clk), .QN(n15449) );
  EDFD1 \Mem_reg[64][0]  ( .D(n24723), .E(n6395), .CP(clk), .QN(n5242) );
  EDFD1 \Mem_reg[63][0]  ( .D(n24723), .E(n6456), .CP(clk), .QN(n5194) );
  EDFD1 \Mem_reg[62][0]  ( .D(n24723), .E(n6455), .CP(clk), .QN(n5146) );
  EDFD1 \Mem_reg[61][0]  ( .D(n24723), .E(n6454), .CP(clk), .QN(n17927) );
  EDFD1 \Mem_reg[60][0]  ( .D(n24723), .E(n6453), .CP(clk), .QN(n17926) );
  EDFD1 \Mem_reg[59][0]  ( .D(n24723), .E(n6452), .CP(clk), .QN(n5002) );
  EDFD1 \Mem_reg[58][0]  ( .D(n24723), .E(n6451), .CP(clk), .QN(n4954) );
  EDFD1 \Mem_reg[57][0]  ( .D(n24723), .E(n6450), .CP(clk), .QN(n4906) );
  EDFD1 \Mem_reg[56][0]  ( .D(n24723), .E(n6449), .CP(clk), .QN(n4858) );
  EDFD1 \Mem_reg[55][0]  ( .D(n24723), .E(n6448), .CP(clk), .QN(n4810) );
  EDFD1 \Mem_reg[54][0]  ( .D(n24723), .E(n6447), .CP(clk), .QN(n15448) );
  EDFD1 \Mem_reg[53][0]  ( .D(n24723), .E(n6446), .CP(clk), .QN(n4714) );
  EDFD1 \Mem_reg[52][0]  ( .D(n24723), .E(n6445), .CP(clk), .Q(n27036) );
  EDFD1 \Mem_reg[51][0]  ( .D(n24723), .E(n6444), .CP(clk), .QN(n4618) );
  EDFD1 \Mem_reg[50][0]  ( .D(n24723), .E(n6443), .CP(clk), .QN(n4570) );
  EDFD1 \Mem_reg[49][0]  ( .D(n24723), .E(n6442), .CP(clk), .QN(n4522) );
  EDFD1 \Mem_reg[48][0]  ( .D(n24723), .E(n6441), .CP(clk), .QN(n4474) );
  EDFD1 \Mem_reg[47][0]  ( .D(n24723), .E(n6440), .CP(clk), .QN(n4426) );
  EDFD1 \Mem_reg[46][0]  ( .D(n24723), .E(n6439), .CP(clk), .QN(n4378) );
  EDFD1 \Mem_reg[43][0]  ( .D(n24723), .E(n6438), .CP(clk), .QN(n4330) );
  EDFD1 \Mem_reg[42][0]  ( .D(n24723), .E(n6437), .CP(clk), .QN(n4282) );
  EDFD1 \Mem_reg[41][0]  ( .D(n24723), .E(n6436), .CP(clk), .QN(n4234) );
  EDFD1 \Mem_reg[40][0]  ( .D(n24723), .E(n6435), .CP(clk), .QN(n4186) );
  EDFD1 \Mem_reg[39][0]  ( .D(n24723), .E(n6434), .CP(clk), .QN(n4138) );
  EDFD1 \Mem_reg[38][0]  ( .D(n24723), .E(n6433), .CP(clk), .QN(n4090) );
  EDFD1 \Mem_reg[37][0]  ( .D(n24723), .E(n6432), .CP(clk), .QN(n4042) );
  EDFD1 \Mem_reg[36][0]  ( .D(n24723), .E(n6431), .CP(clk), .QN(n3994) );
  EDFD1 \Mem_reg[35][0]  ( .D(n24723), .E(n6430), .CP(clk), .QN(n3946) );
  EDFD1 \Mem_reg[34][0]  ( .D(n24723), .E(n6429), .CP(clk), .QN(n3898) );
  EDFD1 \Mem_reg[33][0]  ( .D(n24723), .E(n6428), .CP(clk), .QN(n3850) );
  EDFD1 \Mem_reg[32][0]  ( .D(n24723), .E(n6427), .CP(clk), .QN(n3802) );
  EDFD1 \Mem_reg[31][0]  ( .D(n24723), .E(n6426), .CP(clk), .QN(n3754) );
  EDFD1 \Mem_reg[30][0]  ( .D(n24723), .E(n6425), .CP(clk), .QN(n3706) );
  EDFD1 \Mem_reg[29][0]  ( .D(n24723), .E(n6424), .CP(clk), .QN(n3658) );
  EDFD1 \Mem_reg[28][0]  ( .D(n24723), .E(n6423), .CP(clk), .QN(n3610) );
  EDFD1 \Mem_reg[27][0]  ( .D(n24723), .E(n6422), .CP(clk), .QN(n3562) );
  EDFD1 \Mem_reg[26][0]  ( .D(n24723), .E(n6421), .CP(clk), .QN(n3514) );
  EDFD1 \Mem_reg[25][0]  ( .D(n24723), .E(n6420), .CP(clk), .QN(n3466) );
  EDFD1 \Mem_reg[24][0]  ( .D(n24723), .E(n6463), .CP(clk), .QN(n3418) );
  EDFD1 \Mem_reg[23][0]  ( .D(n24723), .E(n6464), .CP(clk), .QN(n3370) );
  EDFD1 \Mem_reg[22][0]  ( .D(n24723), .E(n6465), .CP(clk), .QN(n3322) );
  EDFD1 \Mem_reg[21][0]  ( .D(n24723), .E(n6466), .CP(clk), .QN(n3274) );
  EDFD1 \Mem_reg[20][0]  ( .D(n24723), .E(n6467), .CP(clk), .QN(n3226) );
  EDFD1 \Mem_reg[19][0]  ( .D(n24723), .E(n6468), .CP(clk), .QN(n3178) );
  EDFD1 \Mem_reg[18][0]  ( .D(n24723), .E(n6469), .CP(clk), .QN(n3130) );
  EDFD1 \Mem_reg[17][0]  ( .D(n24723), .E(n6470), .CP(clk), .QN(n3082) );
  EDFD1 \Mem_reg[16][0]  ( .D(n24723), .E(n6471), .CP(clk), .QN(n3034) );
  EDFD1 \Mem_reg[15][0]  ( .D(n24723), .E(n6472), .CP(clk), .QN(n2986) );
  EDFD1 \Mem_reg[14][0]  ( .D(n24723), .E(n24720), .CP(clk), .QN(n2938) );
  EDFD1 \Mem_reg[13][0]  ( .D(n24723), .E(n24709), .CP(clk), .QN(n2890) );
  EDFD1 \Mem_reg[12][0]  ( .D(n24723), .E(n24717), .CP(clk), .QN(n2842) );
  EDFD1 \Mem_reg[11][0]  ( .D(n24723), .E(n24707), .CP(clk), .QN(n2794) );
  EDFD1 \Mem_reg[10][0]  ( .D(n24723), .E(n6477), .CP(clk), .QN(n2746) );
  EDFD1 \Mem_reg[9][0]  ( .D(n24723), .E(n24708), .CP(clk), .QN(n2698) );
  EDFD1 \Mem_reg[8][0]  ( .D(n24723), .E(n15642), .CP(clk), .QN(n2650) );
  EDFD1 \Mem_reg[7][0]  ( .D(n24723), .E(n24718), .CP(clk), .QN(n2602) );
  EDFD1 \Mem_reg[6][0]  ( .D(n24723), .E(n24716), .CP(clk), .QN(n2554) );
  EDFD1 \Mem_reg[5][0]  ( .D(n24723), .E(n24719), .CP(clk), .QN(n2506) );
  EDFD1 \Mem_reg[4][0]  ( .D(n24723), .E(n24706), .CP(clk), .QN(n2458) );
  EDFD1 \Mem_reg[3][0]  ( .D(n24723), .E(n24721), .CP(clk), .QN(n2410) );
  EDFD1 \Mem_reg[2][0]  ( .D(n24723), .E(n6460), .CP(clk), .QN(n2362) );
  EDFD1 \Mem_reg[1][0]  ( .D(n24723), .E(n24703), .CP(clk), .QN(n2314) );
  EDFD1 \Mem_reg[0][0]  ( .D(n24723), .E(n24705), .CP(clk), .QN(n2266) );
  NR3D0 U7401 ( .A1(Address[5]), .A2(Address[6]), .A3(Address[4]), .ZN(n26975)
         );
  OR2D1 U7402 ( .A1(n24919), .A2(n25068), .Z(n24710) );
  OR2D1 U7403 ( .A1(n24919), .A2(n25070), .Z(n24711) );
  OR2D1 U7404 ( .A1(n24919), .A2(n24920), .Z(n24712) );
  OR2D1 U7405 ( .A1(n24919), .A2(n24965), .Z(n24713) );
  OR2D1 U7406 ( .A1(n24919), .A2(n24922), .Z(n24714) );
  OR2D1 U7407 ( .A1(n24919), .A2(n25069), .Z(n24715) );
  ND2D1 U7408 ( .A1(n26992), .A2(n26975), .ZN(n25068) );
  ND2D1 U7409 ( .A1(n26975), .A2(n26989), .ZN(n24922) );
  CKND0 U7410 ( .I(n24915), .ZN(n26989) );
  ND2D1 U7411 ( .A1(n26975), .A2(n26979), .ZN(n24920) );
  CKND0 U7412 ( .I(n24942), .ZN(n26979) );
  ND2D1 U7413 ( .A1(n26991), .A2(n26975), .ZN(n24965) );
  ND2D1 U7414 ( .A1(n26998), .A2(n26975), .ZN(n25070) );
  ND2D1 U7415 ( .A1(n26983), .A2(n26975), .ZN(n25069) );
  ND2D1 U7416 ( .A1(n26979), .A2(n24952), .ZN(n25063) );
  NR2D2 U7417 ( .A1(n24915), .A2(n24916), .ZN(n24819) );
  NR2D2 U7418 ( .A1(n24918), .A2(n24916), .ZN(n24821) );
  INVD1 U7419 ( .I(n24712), .ZN(n24716) );
  NR2D2 U7420 ( .A1(n24919), .A2(n24921), .ZN(n6477) );
  INVD1 U7421 ( .I(n24714), .ZN(n24717) );
  NR2D2 U7422 ( .A1(n24919), .A2(n24923), .ZN(n6472) );
  NR2D2 U7423 ( .A1(n24919), .A2(n24924), .ZN(n6471) );
  NR2D2 U7424 ( .A1(n24919), .A2(n24925), .ZN(n6470) );
  NR2D2 U7425 ( .A1(n24919), .A2(n24926), .ZN(n6469) );
  NR2D2 U7426 ( .A1(n24919), .A2(n24927), .ZN(n6468) );
  NR2D2 U7427 ( .A1(n24919), .A2(n24928), .ZN(n6467) );
  NR2D2 U7428 ( .A1(n24919), .A2(n24929), .ZN(n6466) );
  NR2D2 U7429 ( .A1(n24919), .A2(n24930), .ZN(n6465) );
  NR2D2 U7430 ( .A1(n24919), .A2(n24931), .ZN(n6464) );
  NR2D2 U7431 ( .A1(n24919), .A2(n24932), .ZN(n6463) );
  NR2D2 U7432 ( .A1(n24919), .A2(n24933), .ZN(n6460) );
  NR2D2 U7433 ( .A1(n24934), .A2(n24935), .ZN(n6456) );
  NR2D2 U7434 ( .A1(n24938), .A2(n24935), .ZN(n6451) );
  NR2D2 U7435 ( .A1(n24940), .A2(n24935), .ZN(n6449) );
  NR2D2 U7436 ( .A1(n24944), .A2(n24935), .ZN(n6445) );
  NR2D2 U7437 ( .A1(n24945), .A2(n24935), .ZN(n6444) );
  NR2D2 U7438 ( .A1(n24946), .A2(n24935), .ZN(n6443) );
  NR2XD1 U7439 ( .A1(n24948), .A2(n24935), .ZN(n6441) );
  ND3D1 U7440 ( .A1(n24949), .A2(n24950), .A3(n24951), .ZN(n24935) );
  NR2D2 U7441 ( .A1(n24916), .A2(n24936), .ZN(n6439) );
  NR2XD1 U7442 ( .A1(n24916), .A2(n24937), .ZN(n6438) );
  ND3D1 U7443 ( .A1(n24952), .A2(n24950), .A3(n24949), .ZN(n24916) );
  NR2D2 U7444 ( .A1(n24916), .A2(n24942), .ZN(n6433) );
  NR2D2 U7445 ( .A1(n24916), .A2(n24943), .ZN(n6432) );
  NR2D2 U7446 ( .A1(n24916), .A2(n24947), .ZN(n6428) );
  NR2D2 U7447 ( .A1(n24934), .A2(n24958), .ZN(n6410) );
  NR2D2 U7448 ( .A1(n24936), .A2(n24958), .ZN(n6409) );
  NR2D2 U7449 ( .A1(n24938), .A2(n24958), .ZN(n6405) );
  NR2D2 U7450 ( .A1(n24939), .A2(n24958), .ZN(n6404) );
  NR2D2 U7451 ( .A1(n24940), .A2(n24958), .ZN(n6403) );
  NR2D2 U7452 ( .A1(n24941), .A2(n24958), .ZN(n6402) );
  NR2D2 U7453 ( .A1(n24919), .A2(n24960), .ZN(n24709) );
  NR2D2 U7454 ( .A1(n24919), .A2(n24961), .ZN(n24708) );
  NR2D2 U7455 ( .A1(n24919), .A2(n24962), .ZN(n24707) );
  NR2D2 U7456 ( .A1(n24919), .A2(n24963), .ZN(n24706) );
  NR2D2 U7457 ( .A1(n24919), .A2(n24964), .ZN(n24705) );
  INVD1 U7458 ( .I(n24713), .ZN(n24718) );
  NR2D2 U7459 ( .A1(n24919), .A2(n24966), .ZN(n24703) );
  INVD1 U7460 ( .I(n24711), .ZN(n24719) );
  NR2D2 U7461 ( .A1(n24919), .A2(n25072), .ZN(n15642) );
  INVD1 U7462 ( .I(n24715), .ZN(n24720) );
  INVD1 U7463 ( .I(n24710), .ZN(n24721) );
  NR2D3 U7464 ( .A1(OE), .A2(CS), .ZN(n2209) );
  CKND0 U7465 ( .I(n15660), .ZN(n24722) );
  INVD1 U7466 ( .I(n24722), .ZN(n24723) );
  CKND0 U7467 ( .I(n15662), .ZN(n24724) );
  INVD1 U7468 ( .I(n24724), .ZN(n24725) );
  CKND0 U7469 ( .I(n15664), .ZN(n24726) );
  INVD1 U7470 ( .I(n24726), .ZN(n24727) );
  CKND0 U7471 ( .I(n15666), .ZN(n24728) );
  INVD1 U7472 ( .I(n24728), .ZN(n24729) );
  CKND0 U7473 ( .I(n15668), .ZN(n24730) );
  INVD1 U7474 ( .I(n24730), .ZN(n24731) );
  CKND0 U7475 ( .I(n15670), .ZN(n24732) );
  INVD1 U7476 ( .I(n24732), .ZN(n24733) );
  CKND0 U7477 ( .I(n15672), .ZN(n24734) );
  INVD1 U7478 ( .I(n24734), .ZN(n24735) );
  CKND0 U7479 ( .I(n15674), .ZN(n24736) );
  INVD1 U7480 ( .I(n24736), .ZN(n24737) );
  CKND0 U7481 ( .I(n15676), .ZN(n24738) );
  INVD1 U7482 ( .I(n24738), .ZN(n24739) );
  CKND0 U7483 ( .I(n15678), .ZN(n24740) );
  INVD1 U7484 ( .I(n24740), .ZN(n24741) );
  CKND0 U7485 ( .I(n15680), .ZN(n24742) );
  INVD1 U7486 ( .I(n24742), .ZN(n24743) );
  CKND0 U7487 ( .I(n15682), .ZN(n24744) );
  INVD1 U7488 ( .I(n24744), .ZN(n24745) );
  CKND0 U7489 ( .I(n15684), .ZN(n24746) );
  INVD1 U7490 ( .I(n24746), .ZN(n24747) );
  CKND0 U7491 ( .I(n15686), .ZN(n24748) );
  INVD1 U7492 ( .I(n24748), .ZN(n24749) );
  CKND0 U7493 ( .I(n15688), .ZN(n24750) );
  INVD1 U7494 ( .I(n24750), .ZN(n24751) );
  CKND0 U7495 ( .I(n15690), .ZN(n24752) );
  INVD1 U7496 ( .I(n24752), .ZN(n24753) );
  CKND0 U7497 ( .I(n15692), .ZN(n24754) );
  INVD1 U7498 ( .I(n24754), .ZN(n24755) );
  CKND0 U7499 ( .I(n15694), .ZN(n24756) );
  INVD1 U7500 ( .I(n24756), .ZN(n24757) );
  CKND0 U7501 ( .I(n15696), .ZN(n24758) );
  INVD1 U7502 ( .I(n24758), .ZN(n24759) );
  CKND0 U7503 ( .I(n15698), .ZN(n24760) );
  INVD1 U7504 ( .I(n24760), .ZN(n24761) );
  CKND0 U7505 ( .I(n15700), .ZN(n24762) );
  INVD1 U7506 ( .I(n24762), .ZN(n24763) );
  CKND0 U7507 ( .I(n15702), .ZN(n24764) );
  INVD1 U7508 ( .I(n24764), .ZN(n24765) );
  CKND0 U7509 ( .I(n15704), .ZN(n24766) );
  INVD1 U7510 ( .I(n24766), .ZN(n24767) );
  CKND0 U7511 ( .I(n15706), .ZN(n24768) );
  INVD1 U7512 ( .I(n24768), .ZN(n24769) );
  CKND0 U7513 ( .I(n15708), .ZN(n24770) );
  INVD1 U7514 ( .I(n24770), .ZN(n24771) );
  CKND0 U7515 ( .I(n15710), .ZN(n24772) );
  INVD1 U7516 ( .I(n24772), .ZN(n24773) );
  CKND0 U7517 ( .I(n15712), .ZN(n24774) );
  INVD1 U7518 ( .I(n24774), .ZN(n24775) );
  CKND0 U7519 ( .I(n15714), .ZN(n24776) );
  INVD1 U7520 ( .I(n24776), .ZN(n24777) );
  CKND0 U7521 ( .I(n15716), .ZN(n24778) );
  INVD1 U7522 ( .I(n24778), .ZN(n24779) );
  CKND0 U7523 ( .I(n15718), .ZN(n24780) );
  INVD1 U7524 ( .I(n24780), .ZN(n24781) );
  CKND0 U7525 ( .I(n15720), .ZN(n24782) );
  INVD1 U7526 ( .I(n24782), .ZN(n24783) );
  CKND0 U7527 ( .I(n15722), .ZN(n24784) );
  INVD1 U7528 ( .I(n24784), .ZN(n24785) );
  CKND0 U7529 ( .I(n15724), .ZN(n24786) );
  INVD1 U7530 ( .I(n24786), .ZN(n24787) );
  CKND0 U7531 ( .I(n15726), .ZN(n24788) );
  INVD1 U7532 ( .I(n24788), .ZN(n24789) );
  CKND0 U7533 ( .I(n15728), .ZN(n24790) );
  INVD1 U7534 ( .I(n24790), .ZN(n24791) );
  CKND0 U7535 ( .I(n15730), .ZN(n24792) );
  INVD1 U7536 ( .I(n24792), .ZN(n24793) );
  CKND0 U7537 ( .I(n15732), .ZN(n24794) );
  INVD1 U7538 ( .I(n24794), .ZN(n24795) );
  CKND0 U7539 ( .I(n15734), .ZN(n24796) );
  INVD1 U7540 ( .I(n24796), .ZN(n24797) );
  CKND0 U7541 ( .I(n15736), .ZN(n24798) );
  INVD1 U7542 ( .I(n24798), .ZN(n24799) );
  CKND0 U7543 ( .I(n15738), .ZN(n24800) );
  INVD1 U7544 ( .I(n24800), .ZN(n24801) );
  CKND0 U7545 ( .I(n15740), .ZN(n24802) );
  INVD1 U7546 ( .I(n24802), .ZN(n24803) );
  CKND0 U7547 ( .I(n15742), .ZN(n24804) );
  INVD1 U7548 ( .I(n24804), .ZN(n24805) );
  CKND0 U7549 ( .I(n15744), .ZN(n24806) );
  INVD1 U7550 ( .I(n24806), .ZN(n24807) );
  CKND0 U7551 ( .I(n15746), .ZN(n24808) );
  INVD1 U7552 ( .I(n24808), .ZN(n24809) );
  CKND0 U7553 ( .I(n15748), .ZN(n24810) );
  INVD1 U7554 ( .I(n24810), .ZN(n24811) );
  CKND0 U7555 ( .I(n15750), .ZN(n24812) );
  INVD1 U7556 ( .I(n24812), .ZN(n24813) );
  CKND0 U7557 ( .I(n15752), .ZN(n24814) );
  INVD1 U7558 ( .I(n24814), .ZN(n24815) );
  CKND0 U7559 ( .I(n15754), .ZN(n24816) );
  INVD1 U7560 ( .I(n24816), .ZN(n24817) );
  ND2D1 U7561 ( .A1(n26976), .A2(n26975), .ZN(n24966) );
  ND2D1 U7562 ( .A1(n26980), .A2(n24951), .ZN(n24984) );
  ND2D1 U7563 ( .A1(n26992), .A2(n24952), .ZN(n25060) );
  NR2D2 U7564 ( .A1(n24942), .A2(n24958), .ZN(n6401) );
  NR2D2 U7565 ( .A1(n24946), .A2(n24955), .ZN(n6413) );
  NR2XD1 U7566 ( .A1(n24937), .A2(n24958), .ZN(n6406) );
  ND3D1 U7567 ( .A1(n24949), .A2(n24956), .A3(n24959), .ZN(n24958) );
  NR2D2 U7568 ( .A1(n24915), .A2(n24935), .ZN(n6453) );
  NR2D2 U7569 ( .A1(n24916), .A2(n24939), .ZN(n6436) );
  ND2D1 U7570 ( .A1(n26977), .A2(n24954), .ZN(n24928) );
  ND2D1 U7571 ( .A1(n24951), .A2(n26990), .ZN(n24994) );
  ND2D1 U7572 ( .A1(n26980), .A2(n24952), .ZN(n25074) );
  ND2D1 U7573 ( .A1(n26982), .A2(n26975), .ZN(n24921) );
  ND2D1 U7574 ( .A1(n27013), .A2(n26975), .ZN(n25072) );
  NR2D2 U7575 ( .A1(n24941), .A2(n24955), .ZN(n6418) );
  NR2D2 U7576 ( .A1(n24944), .A2(n24958), .ZN(n6399) );
  NR2D2 U7577 ( .A1(n24943), .A2(n24935), .ZN(n6446) );
  NR2D2 U7578 ( .A1(n24916), .A2(n24945), .ZN(n6430) );
  ND2D1 U7579 ( .A1(n26983), .A2(n24952), .ZN(n24987) );
  ND2D1 U7580 ( .A1(n24951), .A2(n26998), .ZN(n25048) );
  CKND2D1 U7581 ( .A1(n26977), .A2(n26975), .ZN(n24963) );
  NR2D2 U7582 ( .A1(n24948), .A2(n24955), .ZN(n6411) );
  NR2D2 U7583 ( .A1(n24918), .A2(n24958), .ZN(n6408) );
  NR2D2 U7584 ( .A1(n24938), .A2(n24953), .ZN(n6421) );
  NR2D2 U7585 ( .A1(n24947), .A2(n24935), .ZN(n6442) );
  NR2D2 U7586 ( .A1(n24916), .A2(n24934), .ZN(n6440) );
  ND2D1 U7587 ( .A1(n27013), .A2(n24954), .ZN(n24932) );
  ND2D1 U7588 ( .A1(n24951), .A2(n26979), .ZN(n24997) );
  ND2D1 U7589 ( .A1(n26974), .A2(n26975), .ZN(n24964) );
  ND2D1 U7590 ( .A1(n26989), .A2(n24952), .ZN(n25040) );
  ND2D1 U7591 ( .A1(n26981), .A2(n24951), .ZN(n24983) );
  NR2XD0 U7592 ( .A1(n27023), .A2(n24956), .ZN(n24951) );
  NR2D2 U7593 ( .A1(n24942), .A2(n24955), .ZN(n6417) );
  NR2D2 U7594 ( .A1(n24937), .A2(n24953), .ZN(n6422) );
  NR2D2 U7595 ( .A1(n24915), .A2(n24958), .ZN(n6407) );
  NR2D2 U7596 ( .A1(n24941), .A2(n24935), .ZN(n6448) );
  NR2D2 U7597 ( .A1(n24916), .A2(n24940), .ZN(n6435) );
  ND2D1 U7598 ( .A1(n26992), .A2(n24954), .ZN(n24927) );
  ND2D1 U7599 ( .A1(n24959), .A2(n26977), .ZN(n25024) );
  ND2D1 U7600 ( .A1(n26997), .A2(n26975), .ZN(n24933) );
  ND2D1 U7601 ( .A1(n26990), .A2(n24952), .ZN(n25047) );
  ND2D1 U7602 ( .A1(n24951), .A2(n26974), .ZN(n24980) );
  ND2D1 U7603 ( .A1(n27013), .A2(n24952), .ZN(n25062) );
  NR2XD0 U7604 ( .A1(n24956), .A2(Address[4]), .ZN(n24952) );
  NR2D2 U7605 ( .A1(n24944), .A2(n24955), .ZN(n6415) );
  NR2D2 U7606 ( .A1(n24948), .A2(n24958), .ZN(n6395) );
  NR2D2 U7607 ( .A1(n24939), .A2(n24953), .ZN(n6420) );
  NR2D2 U7608 ( .A1(n24918), .A2(n24935), .ZN(n6454) );
  NR2D2 U7609 ( .A1(n24916), .A2(n24946), .ZN(n6429) );
  ND2D1 U7610 ( .A1(n26976), .A2(n24954), .ZN(n24925) );
  ND2D1 U7611 ( .A1(n26981), .A2(n26988), .ZN(n25005) );
  ND2D1 U7612 ( .A1(n24959), .A2(n26992), .ZN(n25037) );
  ND2D1 U7613 ( .A1(n26975), .A2(n26990), .ZN(n24960) );
  ND2D1 U7614 ( .A1(n26998), .A2(n24952), .ZN(n25059) );
  ND2D1 U7615 ( .A1(n24951), .A2(n26991), .ZN(n24996) );
  CKND0 U7616 ( .I(n24941), .ZN(n26991) );
  NR2D2 U7617 ( .A1(n24943), .A2(n24955), .ZN(n6416) );
  NR2D2 U7618 ( .A1(n24945), .A2(n24958), .ZN(n6398) );
  NR2D2 U7619 ( .A1(n24942), .A2(n24935), .ZN(n6447) );
  NR2D2 U7620 ( .A1(n24934), .A2(n24953), .ZN(n6426) );
  NR2D2 U7621 ( .A1(n24916), .A2(n24938), .ZN(n6437) );
  ND2D1 U7622 ( .A1(n26983), .A2(n26988), .ZN(n25007) );
  ND2D1 U7623 ( .A1(n27003), .A2(n27018), .ZN(n25034) );
  ND2D1 U7624 ( .A1(n24959), .A2(n27013), .ZN(n25027) );
  ND2D1 U7625 ( .A1(n24954), .A2(n26974), .ZN(n24924) );
  ND2D1 U7626 ( .A1(n26981), .A2(n24952), .ZN(n25071) );
  ND2D1 U7627 ( .A1(n24951), .A2(n26997), .ZN(n25036) );
  CKND0 U7628 ( .I(n24946), .ZN(n26997) );
  ND2D1 U7629 ( .A1(n26980), .A2(n26975), .ZN(n24961) );
  NR2D2 U7630 ( .A1(n24947), .A2(n24955), .ZN(n6412) );
  NR2D2 U7631 ( .A1(n24946), .A2(n24958), .ZN(n6397) );
  NR2D2 U7632 ( .A1(n24915), .A2(n24953), .ZN(n6423) );
  NR2D2 U7633 ( .A1(n24935), .A2(n24936), .ZN(n6455) );
  NR2D2 U7634 ( .A1(n24916), .A2(n24941), .ZN(n6434) );
  AN2XD1 U7635 ( .A1(n24957), .A2(Address[3]), .Z(n25044) );
  NR2XD0 U7636 ( .A1(n24950), .A2(n27023), .ZN(n24957) );
  ND2D1 U7637 ( .A1(n26997), .A2(n24954), .ZN(n24926) );
  ND2D1 U7638 ( .A1(Address[6]), .A2(n26981), .ZN(n25039) );
  ND2D1 U7639 ( .A1(n26991), .A2(n24954), .ZN(n24931) );
  AN2XD1 U7640 ( .A1(n26988), .A2(n24950), .Z(n24954) );
  ND2D1 U7641 ( .A1(n26974), .A2(n24952), .ZN(n24986) );
  ND2D1 U7642 ( .A1(n26988), .A2(n26990), .ZN(n25006) );
  ND2D1 U7643 ( .A1(n27003), .A2(n27012), .ZN(n25023) );
  ND2D1 U7644 ( .A1(n24959), .A2(n26991), .ZN(n25014) );
  ND2D1 U7645 ( .A1(n24951), .A2(n27013), .ZN(n25075) );
  INVD1 U7646 ( .I(n24940), .ZN(n27013) );
  ND2D1 U7647 ( .A1(n26978), .A2(n26975), .ZN(n24923) );
  ND2D1 U7648 ( .A1(n26998), .A2(n24954), .ZN(n24929) );
  NR2D2 U7649 ( .A1(n24936), .A2(n24953), .ZN(n6425) );
  NR2D2 U7650 ( .A1(n24940), .A2(n24955), .ZN(n6419) );
  NR2D2 U7651 ( .A1(n24943), .A2(n24958), .ZN(n6400) );
  NR2D2 U7652 ( .A1(n24935), .A2(n24937), .ZN(n6452) );
  NR2D2 U7653 ( .A1(n24916), .A2(n24944), .ZN(n6431) );
  ND2D1 U7654 ( .A1(Address[6]), .A2(n26980), .ZN(n25038) );
  ND2D1 U7655 ( .A1(Address[6]), .A2(n26978), .ZN(n25057) );
  ND2D1 U7656 ( .A1(Address[6]), .A2(n26989), .ZN(n25042) );
  ND2D1 U7657 ( .A1(n27003), .A2(n27004), .ZN(n25017) );
  ND2D1 U7658 ( .A1(n26997), .A2(n24952), .ZN(n25056) );
  ND2D1 U7659 ( .A1(n24957), .A2(n26974), .ZN(n25016) );
  ND2D1 U7660 ( .A1(n26988), .A2(n26982), .ZN(n25004) );
  INVD1 U7661 ( .I(n24938), .ZN(n26982) );
  ND2D1 U7662 ( .A1(n24959), .A2(n26997), .ZN(n25033) );
  ND2D1 U7663 ( .A1(n24951), .A2(n26978), .ZN(n24981) );
  INVD1 U7664 ( .I(n24934), .ZN(n26978) );
  ND2D1 U7665 ( .A1(Address[6]), .A2(n26990), .ZN(n25041) );
  ND2D1 U7666 ( .A1(n27007), .A2(n27012), .ZN(n25026) );
  ND2D1 U7667 ( .A1(n26981), .A2(n26975), .ZN(n24962) );
  ND2D1 U7668 ( .A1(n24954), .A2(n26979), .ZN(n24930) );
  NR2D2 U7669 ( .A1(n24945), .A2(n24955), .ZN(n6414) );
  NR2D2 U7670 ( .A1(n24947), .A2(n24958), .ZN(n6396) );
  NR2D2 U7671 ( .A1(n24918), .A2(n24953), .ZN(n6424) );
  NR2D2 U7672 ( .A1(n24935), .A2(n24939), .ZN(n6450) );
  NR2D2 U7673 ( .A1(n24916), .A2(n24948), .ZN(n6427) );
  MUX2ND0 U7674 ( .I0(n24818), .I1(n24816), .S(n24819), .ZN(n6577) );
  MUX2ND0 U7675 ( .I0(n24820), .I1(n24816), .S(n24821), .ZN(n6576) );
  MUX2ND0 U7676 ( .I0(n24822), .I1(n24814), .S(n24819), .ZN(n6575) );
  MUX2ND0 U7677 ( .I0(n24823), .I1(n24814), .S(n24821), .ZN(n6574) );
  MUX2ND0 U7678 ( .I0(n24824), .I1(n24812), .S(n24819), .ZN(n6573) );
  MUX2ND0 U7679 ( .I0(n24825), .I1(n24812), .S(n24821), .ZN(n6572) );
  MUX2ND0 U7680 ( .I0(n24826), .I1(n24810), .S(n24819), .ZN(n6571) );
  MUX2ND0 U7681 ( .I0(n24827), .I1(n24810), .S(n24821), .ZN(n6570) );
  MUX2ND0 U7682 ( .I0(n24828), .I1(n24808), .S(n24819), .ZN(n6569) );
  MUX2ND0 U7683 ( .I0(n24829), .I1(n24808), .S(n24821), .ZN(n6568) );
  MUX2ND0 U7684 ( .I0(n24830), .I1(n24806), .S(n24819), .ZN(n6567) );
  MUX2ND0 U7685 ( .I0(n24831), .I1(n24806), .S(n24821), .ZN(n6566) );
  MUX2ND0 U7686 ( .I0(n24832), .I1(n24804), .S(n24819), .ZN(n6565) );
  MUX2ND0 U7687 ( .I0(n24833), .I1(n24804), .S(n24821), .ZN(n6564) );
  MUX2ND0 U7688 ( .I0(n24834), .I1(n24802), .S(n24819), .ZN(n6563) );
  MUX2ND0 U7689 ( .I0(n24835), .I1(n24802), .S(n24821), .ZN(n6562) );
  MUX2ND0 U7690 ( .I0(n24836), .I1(n24800), .S(n24819), .ZN(n6561) );
  MUX2ND0 U7691 ( .I0(n24837), .I1(n24800), .S(n24821), .ZN(n6560) );
  MUX2ND0 U7692 ( .I0(n24838), .I1(n24798), .S(n24819), .ZN(n6559) );
  MUX2ND0 U7693 ( .I0(n24839), .I1(n24798), .S(n24821), .ZN(n6558) );
  MUX2ND0 U7694 ( .I0(n24840), .I1(n24796), .S(n24819), .ZN(n6557) );
  MUX2ND0 U7695 ( .I0(n24841), .I1(n24796), .S(n24821), .ZN(n6556) );
  MUX2ND0 U7696 ( .I0(n24842), .I1(n24794), .S(n24819), .ZN(n6555) );
  MUX2ND0 U7697 ( .I0(n24843), .I1(n24794), .S(n24821), .ZN(n6554) );
  MUX2ND0 U7698 ( .I0(n24844), .I1(n24792), .S(n24819), .ZN(n6553) );
  MUX2ND0 U7699 ( .I0(n24845), .I1(n24792), .S(n24821), .ZN(n6552) );
  MUX2ND0 U7700 ( .I0(n24846), .I1(n24790), .S(n24819), .ZN(n6551) );
  MUX2ND0 U7701 ( .I0(n24847), .I1(n24790), .S(n24821), .ZN(n6550) );
  MUX2ND0 U7702 ( .I0(n24848), .I1(n24788), .S(n24819), .ZN(n6549) );
  MUX2ND0 U7703 ( .I0(n24849), .I1(n24788), .S(n24821), .ZN(n6548) );
  MUX2ND0 U7704 ( .I0(n24850), .I1(n24786), .S(n24819), .ZN(n6547) );
  MUX2ND0 U7705 ( .I0(n24851), .I1(n24786), .S(n24821), .ZN(n6546) );
  MUX2ND0 U7706 ( .I0(n24852), .I1(n24784), .S(n24819), .ZN(n6545) );
  MUX2ND0 U7707 ( .I0(n24853), .I1(n24784), .S(n24821), .ZN(n6544) );
  MUX2ND0 U7708 ( .I0(n24854), .I1(n24782), .S(n24819), .ZN(n6543) );
  MUX2ND0 U7709 ( .I0(n24855), .I1(n24782), .S(n24821), .ZN(n6542) );
  MUX2ND0 U7710 ( .I0(n24856), .I1(n24780), .S(n24819), .ZN(n6541) );
  MUX2ND0 U7711 ( .I0(n24857), .I1(n24780), .S(n24821), .ZN(n6540) );
  MUX2ND0 U7712 ( .I0(n24858), .I1(n24778), .S(n24819), .ZN(n6539) );
  MUX2ND0 U7713 ( .I0(n24859), .I1(n24778), .S(n24821), .ZN(n6538) );
  MUX2ND0 U7714 ( .I0(n24860), .I1(n24776), .S(n24819), .ZN(n6537) );
  MUX2ND0 U7715 ( .I0(n24861), .I1(n24776), .S(n24821), .ZN(n6536) );
  MUX2ND0 U7716 ( .I0(n24862), .I1(n24774), .S(n24819), .ZN(n6535) );
  MUX2ND0 U7717 ( .I0(n24863), .I1(n24774), .S(n24821), .ZN(n6534) );
  MUX2ND0 U7718 ( .I0(n24864), .I1(n24772), .S(n24819), .ZN(n6533) );
  MUX2ND0 U7719 ( .I0(n24865), .I1(n24772), .S(n24821), .ZN(n6532) );
  MUX2ND0 U7720 ( .I0(n24866), .I1(n24770), .S(n24819), .ZN(n6531) );
  MUX2ND0 U7721 ( .I0(n24867), .I1(n24770), .S(n24821), .ZN(n6530) );
  MUX2ND0 U7722 ( .I0(n24868), .I1(n24768), .S(n24819), .ZN(n6529) );
  MUX2ND0 U7723 ( .I0(n24869), .I1(n24768), .S(n24821), .ZN(n6528) );
  MUX2ND0 U7724 ( .I0(n24870), .I1(n24766), .S(n24819), .ZN(n6527) );
  MUX2ND0 U7725 ( .I0(n24871), .I1(n24766), .S(n24821), .ZN(n6526) );
  MUX2ND0 U7726 ( .I0(n24872), .I1(n24764), .S(n24819), .ZN(n6525) );
  MUX2ND0 U7727 ( .I0(n24873), .I1(n24764), .S(n24821), .ZN(n6524) );
  MUX2ND0 U7728 ( .I0(n24874), .I1(n24762), .S(n24819), .ZN(n6523) );
  MUX2ND0 U7729 ( .I0(n24875), .I1(n24762), .S(n24821), .ZN(n6522) );
  MUX2ND0 U7730 ( .I0(n24876), .I1(n24760), .S(n24819), .ZN(n6521) );
  MUX2ND0 U7731 ( .I0(n24877), .I1(n24760), .S(n24821), .ZN(n6520) );
  MUX2ND0 U7732 ( .I0(n24878), .I1(n24758), .S(n24819), .ZN(n6519) );
  MUX2ND0 U7733 ( .I0(n24879), .I1(n24758), .S(n24821), .ZN(n6518) );
  MUX2ND0 U7734 ( .I0(n24880), .I1(n24756), .S(n24819), .ZN(n6517) );
  MUX2ND0 U7735 ( .I0(n24881), .I1(n24756), .S(n24821), .ZN(n6516) );
  MUX2ND0 U7736 ( .I0(n24882), .I1(n24754), .S(n24819), .ZN(n6515) );
  MUX2ND0 U7737 ( .I0(n24883), .I1(n24754), .S(n24821), .ZN(n6514) );
  MUX2ND0 U7738 ( .I0(n24884), .I1(n24752), .S(n24819), .ZN(n6513) );
  MUX2ND0 U7739 ( .I0(n24885), .I1(n24752), .S(n24821), .ZN(n6512) );
  MUX2ND0 U7740 ( .I0(n24886), .I1(n24750), .S(n24819), .ZN(n6511) );
  MUX2ND0 U7741 ( .I0(n24887), .I1(n24750), .S(n24821), .ZN(n6510) );
  MUX2ND0 U7742 ( .I0(n24888), .I1(n24748), .S(n24819), .ZN(n6509) );
  MUX2ND0 U7743 ( .I0(n24889), .I1(n24748), .S(n24821), .ZN(n6508) );
  MUX2ND0 U7744 ( .I0(n24890), .I1(n24746), .S(n24819), .ZN(n6507) );
  MUX2ND0 U7745 ( .I0(n24891), .I1(n24746), .S(n24821), .ZN(n6506) );
  MUX2ND0 U7746 ( .I0(n24892), .I1(n24744), .S(n24819), .ZN(n6505) );
  MUX2ND0 U7747 ( .I0(n24893), .I1(n24744), .S(n24821), .ZN(n6504) );
  MUX2ND0 U7748 ( .I0(n24894), .I1(n24742), .S(n24819), .ZN(n6503) );
  MUX2ND0 U7749 ( .I0(n24895), .I1(n24742), .S(n24821), .ZN(n6502) );
  MUX2ND0 U7750 ( .I0(n24896), .I1(n24740), .S(n24819), .ZN(n6501) );
  MUX2ND0 U7751 ( .I0(n24897), .I1(n24740), .S(n24821), .ZN(n6500) );
  MUX2ND0 U7752 ( .I0(n24898), .I1(n24738), .S(n24819), .ZN(n6499) );
  MUX2ND0 U7753 ( .I0(n24899), .I1(n24738), .S(n24821), .ZN(n6498) );
  MUX2ND0 U7754 ( .I0(n24900), .I1(n24736), .S(n24819), .ZN(n6497) );
  MUX2ND0 U7755 ( .I0(n24901), .I1(n24736), .S(n24821), .ZN(n6496) );
  MUX2ND0 U7756 ( .I0(n24902), .I1(n24734), .S(n24819), .ZN(n6495) );
  MUX2ND0 U7757 ( .I0(n24903), .I1(n24734), .S(n24821), .ZN(n6494) );
  MUX2ND0 U7758 ( .I0(n24904), .I1(n24732), .S(n24819), .ZN(n6493) );
  MUX2ND0 U7759 ( .I0(n24905), .I1(n24732), .S(n24821), .ZN(n6492) );
  MUX2ND0 U7760 ( .I0(n24906), .I1(n24730), .S(n24819), .ZN(n6491) );
  MUX2ND0 U7761 ( .I0(n24907), .I1(n24730), .S(n24821), .ZN(n6490) );
  MUX2ND0 U7762 ( .I0(n24908), .I1(n24728), .S(n24819), .ZN(n6489) );
  MUX2ND0 U7763 ( .I0(n24909), .I1(n24728), .S(n24821), .ZN(n6488) );
  MUX2ND0 U7764 ( .I0(n24910), .I1(n24726), .S(n24819), .ZN(n6487) );
  MUX2ND0 U7765 ( .I0(n24911), .I1(n24726), .S(n24821), .ZN(n6486) );
  MUX2ND0 U7766 ( .I0(n24912), .I1(n24724), .S(n24819), .ZN(n6485) );
  MUX2ND0 U7767 ( .I0(n24913), .I1(n24724), .S(n24821), .ZN(n6484) );
  MUX2ND0 U7768 ( .I0(n24914), .I1(n24722), .S(n24819), .ZN(n6483) );
  MUX2ND0 U7769 ( .I0(n24917), .I1(n24722), .S(n24821), .ZN(n6482) );
  CKND2D0 U7770 ( .A1(n24954), .A2(n24949), .ZN(n24953) );
  ND3D0 U7771 ( .A1(n24949), .A2(n24956), .A3(n24957), .ZN(n24955) );
  ND4D0 U7772 ( .A1(n24967), .A2(n24968), .A3(n24969), .A4(n24970), .ZN(n2218)
         );
  AN4D0 U7773 ( .A1(n24971), .A2(n24972), .A3(n24973), .A4(n24974), .Z(n24970)
         );
  NR4D0 U7774 ( .A1(n24975), .A2(n24976), .A3(n24977), .A4(n24978), .ZN(n24974) );
  OAI222D0 U7775 ( .A1(n24979), .A2(n15449), .B1(n24980), .B2(n4474), .C1(
        n24964), .C2(n2266), .ZN(n24978) );
  OAI222D0 U7776 ( .A1(n24920), .A2(n2554), .B1(n24981), .B2(n5194), .C1(
        n24963), .C2(n2458), .ZN(n24977) );
  OAI222D0 U7777 ( .A1(n24982), .A2(n4954), .B1(n24983), .B2(n5002), .C1(
        n24984), .C2(n4906), .ZN(n24976) );
  OAI222D0 U7778 ( .A1(n24985), .A2(n4426), .B1(n24986), .B2(n3802), .C1(
        n24987), .C2(n4378), .ZN(n24975) );
  NR4D0 U7779 ( .A1(n24988), .A2(n24989), .A3(n24990), .A4(n24991), .ZN(n24973) );
  OAI22D0 U7780 ( .A1(n24922), .A2(n2842), .B1(n24992), .B2(n3754), .ZN(n24991) );
  OAI222D0 U7781 ( .A1(n24993), .A2(n17926), .B1(n24962), .B2(n2794), .C1(
        n24994), .C2(n17927), .ZN(n24990) );
  OAI222D0 U7782 ( .A1(n24995), .A2(n5242), .B1(n24961), .B2(n2698), .C1(
        n24921), .C2(n2746), .ZN(n24989) );
  OAI222D0 U7783 ( .A1(n24927), .A2(n3178), .B1(n24996), .B2(n4810), .C1(
        n24997), .C2(n15448), .ZN(n24988) );
  NR4D0 U7784 ( .A1(n24998), .A2(n24999), .A3(n25000), .A4(n25001), .ZN(n24972) );
  OAI22D0 U7785 ( .A1(n24928), .A2(n3226), .B1(n24926), .B2(n3130), .ZN(n25001) );
  OAI222D0 U7786 ( .A1(n25002), .A2(n3466), .B1(n24929), .B2(n3274), .C1(
        n24933), .C2(n2362), .ZN(n25000) );
  OAI222D0 U7787 ( .A1(n25003), .A2(n3610), .B1(n25004), .B2(n3514), .C1(
        n25005), .C2(n3562), .ZN(n24999) );
  OAI222D0 U7788 ( .A1(n24965), .A2(n2602), .B1(n25006), .B2(n3658), .C1(
        n25007), .C2(n3706), .ZN(n24998) );
  NR4D0 U7789 ( .A1(n25008), .A2(n25009), .A3(n25010), .A4(n25011), .ZN(n24971) );
  OAI22D0 U7790 ( .A1(n25012), .A2(n5146), .B1(n24966), .B2(n2314), .ZN(n25011) );
  OAI222D0 U7791 ( .A1(n24925), .A2(n3082), .B1(n24923), .B2(n2986), .C1(
        n24960), .C2(n2890), .ZN(n25010) );
  OAI222D0 U7792 ( .A1(n25013), .A2(n5530), .B1(n25014), .B2(n5578), .C1(
        n24924), .C2(n3034), .ZN(n25009) );
  OAI222D0 U7793 ( .A1(n25015), .A2(n6106), .B1(n25016), .B2(n6010), .C1(
        n25017), .C2(n6154), .ZN(n25008) );
  INR4D0 U7794 ( .A1(n25018), .B1(n25019), .B2(n25020), .B3(n25021), .ZN(
        n24969) );
  OAI222D0 U7795 ( .A1(n25022), .A2(n5482), .B1(n25023), .B2(n6346), .C1(
        n25024), .C2(n5434), .ZN(n25021) );
  OAI222D0 U7796 ( .A1(n25025), .A2(n4522), .B1(n25026), .B2(n24559), .C1(
        n25027), .C2(n5626), .ZN(n25020) );
  OR4D0 U7797 ( .A1(n25028), .A2(n25029), .A3(n25030), .A4(n25031), .Z(n25019)
         );
  OAI222D0 U7798 ( .A1(n25032), .A2(n4618), .B1(n25033), .B2(n5338), .C1(
        n25034), .C2(n6250), .ZN(n25031) );
  OAI222D0 U7799 ( .A1(n25035), .A2(n6202), .B1(n25036), .B2(n4570), .C1(
        n25037), .C2(n5386), .ZN(n25030) );
  OAI22D0 U7800 ( .A1(n27039), .A2(n25038), .B1(n27038), .B2(n25039), .ZN(
        n25029) );
  OAI222D0 U7801 ( .A1(n24914), .A2(n25040), .B1(n25041), .B2(n5866), .C1(
        n25042), .C2(n5818), .ZN(n25028) );
  CKND0 U7802 ( .I(\Mem[44][0] ), .ZN(n24914) );
  AOI221D0 U7803 ( .A1(n27036), .A2(n25043), .B1(n27037), .B2(n25044), .C(
        n25045), .ZN(n25018) );
  OAI222D0 U7804 ( .A1(n25046), .A2(n6058), .B1(n24917), .B2(n25047), .C1(
        n25048), .C2(n4714), .ZN(n25045) );
  CKND0 U7805 ( .I(\Mem[45][0] ), .ZN(n24917) );
  NR4D0 U7806 ( .A1(n25049), .A2(n25050), .A3(n25051), .A4(n25052), .ZN(n24968) );
  OAI22D0 U7807 ( .A1(n25053), .A2(n5914), .B1(n25054), .B2(n5722), .ZN(n25052) );
  OAI222D0 U7808 ( .A1(n25055), .A2(n3850), .B1(n25056), .B2(n3898), .C1(
        n25057), .C2(n5962), .ZN(n25051) );
  OAI222D0 U7809 ( .A1(n25058), .A2(n3994), .B1(n25059), .B2(n4042), .C1(
        n25060), .C2(n3946), .ZN(n25050) );
  OAI222D0 U7810 ( .A1(n25061), .A2(n4138), .B1(n25062), .B2(n4186), .C1(
        n25063), .C2(n4090), .ZN(n25049) );
  NR4D0 U7811 ( .A1(n25064), .A2(n25065), .A3(n25066), .A4(n25067), .ZN(n24967) );
  OAI22D0 U7812 ( .A1(n25068), .A2(n2410), .B1(n25069), .B2(n2938), .ZN(n25067) );
  OAI222D0 U7813 ( .A1(n25070), .A2(n2506), .B1(n25071), .B2(n4330), .C1(
        n25072), .C2(n2650), .ZN(n25066) );
  OAI222D0 U7814 ( .A1(n25073), .A2(n4282), .B1(n24930), .B2(n3322), .C1(
        n25074), .C2(n4234), .ZN(n25065) );
  OAI222D0 U7815 ( .A1(n24932), .A2(n3418), .B1(n25075), .B2(n4858), .C1(
        n24931), .C2(n3370), .ZN(n25064) );
  ND4D0 U7816 ( .A1(n25076), .A2(n25077), .A3(n25078), .A4(n25079), .ZN(n2217)
         );
  AN4D0 U7817 ( .A1(n25080), .A2(n25081), .A3(n25082), .A4(n25083), .Z(n25079)
         );
  NR4D0 U7818 ( .A1(n25084), .A2(n25085), .A3(n25086), .A4(n25087), .ZN(n25083) );
  OAI222D0 U7819 ( .A1(n24979), .A2(n15453), .B1(n24980), .B2(n4473), .C1(
        n24964), .C2(n2265), .ZN(n25087) );
  OAI222D0 U7820 ( .A1(n24920), .A2(n2553), .B1(n24981), .B2(n5193), .C1(
        n24963), .C2(n2457), .ZN(n25086) );
  OAI222D0 U7821 ( .A1(n24982), .A2(n4953), .B1(n24983), .B2(n5001), .C1(
        n24984), .C2(n4905), .ZN(n25085) );
  OAI222D0 U7822 ( .A1(n24985), .A2(n4425), .B1(n24986), .B2(n3801), .C1(
        n24987), .C2(n4377), .ZN(n25084) );
  NR4D0 U7823 ( .A1(n25088), .A2(n25089), .A3(n25090), .A4(n25091), .ZN(n25082) );
  OAI22D0 U7824 ( .A1(n24922), .A2(n2841), .B1(n24992), .B2(n3753), .ZN(n25091) );
  OAI222D0 U7825 ( .A1(n24993), .A2(n17929), .B1(n24962), .B2(n2793), .C1(
        n24994), .C2(n17930), .ZN(n25090) );
  OAI222D0 U7826 ( .A1(n24995), .A2(n5241), .B1(n24961), .B2(n2697), .C1(
        n24921), .C2(n2745), .ZN(n25089) );
  OAI222D0 U7827 ( .A1(n24927), .A2(n3177), .B1(n24996), .B2(n4809), .C1(
        n24997), .C2(n15452), .ZN(n25088) );
  NR4D0 U7828 ( .A1(n25092), .A2(n25093), .A3(n25094), .A4(n25095), .ZN(n25081) );
  OAI22D0 U7829 ( .A1(n24928), .A2(n3225), .B1(n24926), .B2(n3129), .ZN(n25095) );
  OAI222D0 U7830 ( .A1(n25002), .A2(n3465), .B1(n24929), .B2(n3273), .C1(
        n24933), .C2(n2361), .ZN(n25094) );
  OAI222D0 U7831 ( .A1(n25003), .A2(n3609), .B1(n25004), .B2(n3513), .C1(
        n25005), .C2(n3561), .ZN(n25093) );
  OAI222D0 U7832 ( .A1(n24965), .A2(n2601), .B1(n25006), .B2(n3657), .C1(
        n25007), .C2(n3705), .ZN(n25092) );
  NR4D0 U7833 ( .A1(n25096), .A2(n25097), .A3(n25098), .A4(n25099), .ZN(n25080) );
  OAI22D0 U7834 ( .A1(n25012), .A2(n5145), .B1(n24966), .B2(n2313), .ZN(n25099) );
  OAI222D0 U7835 ( .A1(n24925), .A2(n3081), .B1(n24923), .B2(n2985), .C1(
        n24960), .C2(n2889), .ZN(n25098) );
  OAI222D0 U7836 ( .A1(n25013), .A2(n5529), .B1(n25014), .B2(n5577), .C1(
        n24924), .C2(n3033), .ZN(n25097) );
  OAI222D0 U7837 ( .A1(n25015), .A2(n6105), .B1(n25016), .B2(n6009), .C1(
        n25017), .C2(n6153), .ZN(n25096) );
  INR4D0 U7838 ( .A1(n25100), .B1(n25101), .B2(n25102), .B3(n25103), .ZN(
        n25078) );
  OAI222D0 U7839 ( .A1(n25022), .A2(n5481), .B1(n25023), .B2(n6345), .C1(
        n25024), .C2(n5433), .ZN(n25103) );
  OAI222D0 U7840 ( .A1(n25025), .A2(n4521), .B1(n25026), .B2(n24562), .C1(
        n25027), .C2(n5625), .ZN(n25102) );
  OR4D0 U7841 ( .A1(n25104), .A2(n25105), .A3(n25106), .A4(n25107), .Z(n25101)
         );
  OAI222D0 U7842 ( .A1(n25032), .A2(n4617), .B1(n25033), .B2(n5337), .C1(
        n25034), .C2(n6249), .ZN(n25107) );
  OAI222D0 U7843 ( .A1(n25035), .A2(n6201), .B1(n25036), .B2(n4569), .C1(
        n25037), .C2(n5385), .ZN(n25106) );
  OAI22D0 U7844 ( .A1(n27043), .A2(n25038), .B1(n27042), .B2(n25039), .ZN(
        n25105) );
  OAI222D0 U7845 ( .A1(n24912), .A2(n25040), .B1(n25041), .B2(n5865), .C1(
        n25042), .C2(n5817), .ZN(n25104) );
  CKND0 U7846 ( .I(\Mem[44][1] ), .ZN(n24912) );
  AOI221D0 U7847 ( .A1(n27040), .A2(n25043), .B1(n27041), .B2(n25044), .C(
        n25108), .ZN(n25100) );
  OAI222D0 U7848 ( .A1(n25046), .A2(n6057), .B1(n24913), .B2(n25047), .C1(
        n25048), .C2(n4713), .ZN(n25108) );
  CKND0 U7849 ( .I(\Mem[45][1] ), .ZN(n24913) );
  NR4D0 U7850 ( .A1(n25109), .A2(n25110), .A3(n25111), .A4(n25112), .ZN(n25077) );
  OAI22D0 U7851 ( .A1(n25053), .A2(n5913), .B1(n25054), .B2(n5721), .ZN(n25112) );
  OAI222D0 U7852 ( .A1(n25055), .A2(n3849), .B1(n25056), .B2(n3897), .C1(
        n25057), .C2(n5961), .ZN(n25111) );
  OAI222D0 U7853 ( .A1(n25058), .A2(n3993), .B1(n25059), .B2(n4041), .C1(
        n25060), .C2(n3945), .ZN(n25110) );
  OAI222D0 U7854 ( .A1(n25061), .A2(n4137), .B1(n25062), .B2(n4185), .C1(
        n25063), .C2(n4089), .ZN(n25109) );
  NR4D0 U7855 ( .A1(n25113), .A2(n25114), .A3(n25115), .A4(n25116), .ZN(n25076) );
  OAI22D0 U7856 ( .A1(n25068), .A2(n2409), .B1(n25069), .B2(n2937), .ZN(n25116) );
  OAI222D0 U7857 ( .A1(n25070), .A2(n2505), .B1(n25071), .B2(n4329), .C1(
        n25072), .C2(n2649), .ZN(n25115) );
  OAI222D0 U7858 ( .A1(n25073), .A2(n4281), .B1(n24930), .B2(n3321), .C1(
        n25074), .C2(n4233), .ZN(n25114) );
  OAI222D0 U7859 ( .A1(n24932), .A2(n3417), .B1(n25075), .B2(n4857), .C1(
        n24931), .C2(n3369), .ZN(n25113) );
  ND4D0 U7860 ( .A1(n25117), .A2(n25118), .A3(n25119), .A4(n25120), .ZN(n2216)
         );
  AN4D0 U7861 ( .A1(n25121), .A2(n25122), .A3(n25123), .A4(n25124), .Z(n25120)
         );
  NR4D0 U7862 ( .A1(n25125), .A2(n25126), .A3(n25127), .A4(n25128), .ZN(n25124) );
  OAI222D0 U7863 ( .A1(n24979), .A2(n15457), .B1(n24980), .B2(n4472), .C1(
        n24964), .C2(n2264), .ZN(n25128) );
  OAI222D0 U7864 ( .A1(n24920), .A2(n2552), .B1(n24981), .B2(n5192), .C1(
        n24963), .C2(n2456), .ZN(n25127) );
  OAI222D0 U7865 ( .A1(n24982), .A2(n4952), .B1(n24983), .B2(n5000), .C1(
        n24984), .C2(n4904), .ZN(n25126) );
  OAI222D0 U7866 ( .A1(n24985), .A2(n4424), .B1(n24986), .B2(n3800), .C1(
        n24987), .C2(n4376), .ZN(n25125) );
  NR4D0 U7867 ( .A1(n25129), .A2(n25130), .A3(n25131), .A4(n25132), .ZN(n25123) );
  OAI22D0 U7868 ( .A1(n24922), .A2(n2840), .B1(n24992), .B2(n3752), .ZN(n25132) );
  OAI222D0 U7869 ( .A1(n24993), .A2(n17932), .B1(n24962), .B2(n2792), .C1(
        n24994), .C2(n17933), .ZN(n25131) );
  OAI222D0 U7870 ( .A1(n24995), .A2(n5240), .B1(n24961), .B2(n2696), .C1(
        n24921), .C2(n2744), .ZN(n25130) );
  OAI222D0 U7871 ( .A1(n24927), .A2(n3176), .B1(n24996), .B2(n4808), .C1(
        n24997), .C2(n15456), .ZN(n25129) );
  NR4D0 U7872 ( .A1(n25133), .A2(n25134), .A3(n25135), .A4(n25136), .ZN(n25122) );
  OAI22D0 U7873 ( .A1(n24928), .A2(n3224), .B1(n24926), .B2(n3128), .ZN(n25136) );
  OAI222D0 U7874 ( .A1(n25002), .A2(n3464), .B1(n24929), .B2(n3272), .C1(
        n24933), .C2(n2360), .ZN(n25135) );
  OAI222D0 U7875 ( .A1(n25003), .A2(n3608), .B1(n25004), .B2(n3512), .C1(
        n25005), .C2(n3560), .ZN(n25134) );
  OAI222D0 U7876 ( .A1(n24965), .A2(n2600), .B1(n25006), .B2(n3656), .C1(
        n25007), .C2(n3704), .ZN(n25133) );
  NR4D0 U7877 ( .A1(n25137), .A2(n25138), .A3(n25139), .A4(n25140), .ZN(n25121) );
  OAI22D0 U7878 ( .A1(n25012), .A2(n5144), .B1(n24966), .B2(n2312), .ZN(n25140) );
  OAI222D0 U7879 ( .A1(n24925), .A2(n3080), .B1(n24923), .B2(n2984), .C1(
        n24960), .C2(n2888), .ZN(n25139) );
  OAI222D0 U7880 ( .A1(n25013), .A2(n5528), .B1(n25014), .B2(n5576), .C1(
        n24924), .C2(n3032), .ZN(n25138) );
  OAI222D0 U7881 ( .A1(n25015), .A2(n6104), .B1(n25016), .B2(n6008), .C1(
        n25017), .C2(n6152), .ZN(n25137) );
  INR4D0 U7882 ( .A1(n25141), .B1(n25142), .B2(n25143), .B3(n25144), .ZN(
        n25119) );
  OAI222D0 U7883 ( .A1(n25022), .A2(n5480), .B1(n25023), .B2(n6344), .C1(
        n25024), .C2(n5432), .ZN(n25144) );
  OAI222D0 U7884 ( .A1(n25025), .A2(n4520), .B1(n25026), .B2(n24565), .C1(
        n25027), .C2(n5624), .ZN(n25143) );
  OR4D0 U7885 ( .A1(n25145), .A2(n25146), .A3(n25147), .A4(n25148), .Z(n25142)
         );
  OAI222D0 U7886 ( .A1(n25032), .A2(n4616), .B1(n25033), .B2(n5336), .C1(
        n25034), .C2(n6248), .ZN(n25148) );
  OAI222D0 U7887 ( .A1(n25035), .A2(n6200), .B1(n25036), .B2(n4568), .C1(
        n25037), .C2(n5384), .ZN(n25147) );
  OAI22D0 U7888 ( .A1(n27047), .A2(n25038), .B1(n27046), .B2(n25039), .ZN(
        n25146) );
  OAI222D0 U7889 ( .A1(n24910), .A2(n25040), .B1(n25041), .B2(n5864), .C1(
        n25042), .C2(n5816), .ZN(n25145) );
  CKND0 U7890 ( .I(\Mem[44][2] ), .ZN(n24910) );
  AOI221D0 U7891 ( .A1(n27044), .A2(n25043), .B1(n27045), .B2(n25044), .C(
        n25149), .ZN(n25141) );
  OAI222D0 U7892 ( .A1(n25046), .A2(n6056), .B1(n24911), .B2(n25047), .C1(
        n25048), .C2(n4712), .ZN(n25149) );
  CKND0 U7893 ( .I(\Mem[45][2] ), .ZN(n24911) );
  NR4D0 U7894 ( .A1(n25150), .A2(n25151), .A3(n25152), .A4(n25153), .ZN(n25118) );
  OAI22D0 U7895 ( .A1(n25053), .A2(n5912), .B1(n25054), .B2(n5720), .ZN(n25153) );
  OAI222D0 U7896 ( .A1(n25055), .A2(n3848), .B1(n25056), .B2(n3896), .C1(
        n25057), .C2(n5960), .ZN(n25152) );
  OAI222D0 U7897 ( .A1(n25058), .A2(n3992), .B1(n25059), .B2(n4040), .C1(
        n25060), .C2(n3944), .ZN(n25151) );
  OAI222D0 U7898 ( .A1(n25061), .A2(n4136), .B1(n25062), .B2(n4184), .C1(
        n25063), .C2(n4088), .ZN(n25150) );
  NR4D0 U7899 ( .A1(n25154), .A2(n25155), .A3(n25156), .A4(n25157), .ZN(n25117) );
  OAI22D0 U7900 ( .A1(n25068), .A2(n2408), .B1(n25069), .B2(n2936), .ZN(n25157) );
  OAI222D0 U7901 ( .A1(n25070), .A2(n2504), .B1(n25071), .B2(n4328), .C1(
        n25072), .C2(n2648), .ZN(n25156) );
  OAI222D0 U7902 ( .A1(n25073), .A2(n4280), .B1(n24930), .B2(n3320), .C1(
        n25074), .C2(n4232), .ZN(n25155) );
  OAI222D0 U7903 ( .A1(n24932), .A2(n3416), .B1(n25075), .B2(n4856), .C1(
        n24931), .C2(n3368), .ZN(n25154) );
  ND4D0 U7904 ( .A1(n25158), .A2(n25159), .A3(n25160), .A4(n25161), .ZN(n2215)
         );
  AN4D0 U7905 ( .A1(n25162), .A2(n25163), .A3(n25164), .A4(n25165), .Z(n25161)
         );
  NR4D0 U7906 ( .A1(n25166), .A2(n25167), .A3(n25168), .A4(n25169), .ZN(n25165) );
  OAI222D0 U7907 ( .A1(n24979), .A2(n15461), .B1(n24980), .B2(n4471), .C1(
        n24964), .C2(n2263), .ZN(n25169) );
  OAI222D0 U7908 ( .A1(n24920), .A2(n2551), .B1(n24981), .B2(n5191), .C1(
        n24963), .C2(n2455), .ZN(n25168) );
  OAI222D0 U7909 ( .A1(n24982), .A2(n4951), .B1(n24983), .B2(n4999), .C1(
        n24984), .C2(n4903), .ZN(n25167) );
  OAI222D0 U7910 ( .A1(n24985), .A2(n4423), .B1(n24986), .B2(n3799), .C1(
        n24987), .C2(n4375), .ZN(n25166) );
  NR4D0 U7911 ( .A1(n25170), .A2(n25171), .A3(n25172), .A4(n25173), .ZN(n25164) );
  OAI22D0 U7912 ( .A1(n24922), .A2(n2839), .B1(n24992), .B2(n3751), .ZN(n25173) );
  OAI222D0 U7913 ( .A1(n24993), .A2(n17935), .B1(n24962), .B2(n2791), .C1(
        n24994), .C2(n17936), .ZN(n25172) );
  OAI222D0 U7914 ( .A1(n24995), .A2(n5239), .B1(n24961), .B2(n2695), .C1(
        n24921), .C2(n2743), .ZN(n25171) );
  OAI222D0 U7915 ( .A1(n24927), .A2(n3175), .B1(n24996), .B2(n4807), .C1(
        n24997), .C2(n15460), .ZN(n25170) );
  NR4D0 U7916 ( .A1(n25174), .A2(n25175), .A3(n25176), .A4(n25177), .ZN(n25163) );
  OAI22D0 U7917 ( .A1(n24928), .A2(n3223), .B1(n24926), .B2(n3127), .ZN(n25177) );
  OAI222D0 U7918 ( .A1(n25002), .A2(n3463), .B1(n24929), .B2(n3271), .C1(
        n24933), .C2(n2359), .ZN(n25176) );
  OAI222D0 U7919 ( .A1(n25003), .A2(n3607), .B1(n25004), .B2(n3511), .C1(
        n25005), .C2(n3559), .ZN(n25175) );
  OAI222D0 U7920 ( .A1(n24965), .A2(n2599), .B1(n25006), .B2(n3655), .C1(
        n25007), .C2(n3703), .ZN(n25174) );
  NR4D0 U7921 ( .A1(n25178), .A2(n25179), .A3(n25180), .A4(n25181), .ZN(n25162) );
  OAI22D0 U7922 ( .A1(n25012), .A2(n5143), .B1(n24966), .B2(n2311), .ZN(n25181) );
  OAI222D0 U7923 ( .A1(n24925), .A2(n3079), .B1(n24923), .B2(n2983), .C1(
        n24960), .C2(n2887), .ZN(n25180) );
  OAI222D0 U7924 ( .A1(n25013), .A2(n5527), .B1(n25014), .B2(n5575), .C1(
        n24924), .C2(n3031), .ZN(n25179) );
  OAI222D0 U7925 ( .A1(n25015), .A2(n6103), .B1(n25016), .B2(n6007), .C1(
        n25017), .C2(n6151), .ZN(n25178) );
  INR4D0 U7926 ( .A1(n25182), .B1(n25183), .B2(n25184), .B3(n25185), .ZN(
        n25160) );
  OAI222D0 U7927 ( .A1(n25022), .A2(n5479), .B1(n25023), .B2(n6343), .C1(
        n25024), .C2(n5431), .ZN(n25185) );
  OAI222D0 U7928 ( .A1(n25025), .A2(n4519), .B1(n25026), .B2(n24568), .C1(
        n25027), .C2(n5623), .ZN(n25184) );
  OR4D0 U7929 ( .A1(n25186), .A2(n25187), .A3(n25188), .A4(n25189), .Z(n25183)
         );
  OAI222D0 U7930 ( .A1(n25032), .A2(n4615), .B1(n25033), .B2(n5335), .C1(
        n25034), .C2(n6247), .ZN(n25189) );
  OAI222D0 U7931 ( .A1(n25035), .A2(n6199), .B1(n25036), .B2(n4567), .C1(
        n25037), .C2(n5383), .ZN(n25188) );
  OAI22D0 U7932 ( .A1(n27051), .A2(n25038), .B1(n27050), .B2(n25039), .ZN(
        n25187) );
  OAI222D0 U7933 ( .A1(n24908), .A2(n25040), .B1(n25041), .B2(n5863), .C1(
        n25042), .C2(n5815), .ZN(n25186) );
  CKND0 U7934 ( .I(\Mem[44][3] ), .ZN(n24908) );
  AOI221D0 U7935 ( .A1(n27048), .A2(n25043), .B1(n27049), .B2(n25044), .C(
        n25190), .ZN(n25182) );
  OAI222D0 U7936 ( .A1(n25046), .A2(n6055), .B1(n24909), .B2(n25047), .C1(
        n25048), .C2(n4711), .ZN(n25190) );
  CKND0 U7937 ( .I(\Mem[45][3] ), .ZN(n24909) );
  NR4D0 U7938 ( .A1(n25191), .A2(n25192), .A3(n25193), .A4(n25194), .ZN(n25159) );
  OAI22D0 U7939 ( .A1(n25053), .A2(n5911), .B1(n25054), .B2(n5719), .ZN(n25194) );
  OAI222D0 U7940 ( .A1(n25055), .A2(n3847), .B1(n25056), .B2(n3895), .C1(
        n25057), .C2(n5959), .ZN(n25193) );
  OAI222D0 U7941 ( .A1(n25058), .A2(n3991), .B1(n25059), .B2(n4039), .C1(
        n25060), .C2(n3943), .ZN(n25192) );
  OAI222D0 U7942 ( .A1(n25061), .A2(n4135), .B1(n25062), .B2(n4183), .C1(
        n25063), .C2(n4087), .ZN(n25191) );
  NR4D0 U7943 ( .A1(n25195), .A2(n25196), .A3(n25197), .A4(n25198), .ZN(n25158) );
  OAI22D0 U7944 ( .A1(n25068), .A2(n2407), .B1(n25069), .B2(n2935), .ZN(n25198) );
  OAI222D0 U7945 ( .A1(n25070), .A2(n2503), .B1(n25071), .B2(n4327), .C1(
        n25072), .C2(n2647), .ZN(n25197) );
  OAI222D0 U7946 ( .A1(n25073), .A2(n4279), .B1(n24930), .B2(n3319), .C1(
        n25074), .C2(n4231), .ZN(n25196) );
  OAI222D0 U7947 ( .A1(n24932), .A2(n3415), .B1(n25075), .B2(n4855), .C1(
        n24931), .C2(n3367), .ZN(n25195) );
  ND4D0 U7948 ( .A1(n25199), .A2(n25200), .A3(n25201), .A4(n25202), .ZN(n2214)
         );
  AN4D0 U7949 ( .A1(n25203), .A2(n25204), .A3(n25205), .A4(n25206), .Z(n25202)
         );
  NR4D0 U7950 ( .A1(n25207), .A2(n25208), .A3(n25209), .A4(n25210), .ZN(n25206) );
  OAI222D0 U7951 ( .A1(n24979), .A2(n15465), .B1(n24980), .B2(n4470), .C1(
        n24964), .C2(n2262), .ZN(n25210) );
  OAI222D0 U7952 ( .A1(n24920), .A2(n2550), .B1(n24981), .B2(n5190), .C1(
        n24963), .C2(n2454), .ZN(n25209) );
  OAI222D0 U7953 ( .A1(n24982), .A2(n4950), .B1(n24983), .B2(n4998), .C1(
        n24984), .C2(n4902), .ZN(n25208) );
  OAI222D0 U7954 ( .A1(n24985), .A2(n4422), .B1(n24986), .B2(n3798), .C1(
        n24987), .C2(n4374), .ZN(n25207) );
  NR4D0 U7955 ( .A1(n25211), .A2(n25212), .A3(n25213), .A4(n25214), .ZN(n25205) );
  OAI22D0 U7956 ( .A1(n24922), .A2(n2838), .B1(n24992), .B2(n3750), .ZN(n25214) );
  OAI222D0 U7957 ( .A1(n24993), .A2(n17938), .B1(n24962), .B2(n2790), .C1(
        n24994), .C2(n17939), .ZN(n25213) );
  OAI222D0 U7958 ( .A1(n24995), .A2(n5238), .B1(n24961), .B2(n2694), .C1(
        n24921), .C2(n2742), .ZN(n25212) );
  OAI222D0 U7959 ( .A1(n24927), .A2(n3174), .B1(n24996), .B2(n4806), .C1(
        n24997), .C2(n15464), .ZN(n25211) );
  NR4D0 U7960 ( .A1(n25215), .A2(n25216), .A3(n25217), .A4(n25218), .ZN(n25204) );
  OAI22D0 U7961 ( .A1(n24928), .A2(n3222), .B1(n24926), .B2(n3126), .ZN(n25218) );
  OAI222D0 U7962 ( .A1(n25002), .A2(n3462), .B1(n24929), .B2(n3270), .C1(
        n24933), .C2(n2358), .ZN(n25217) );
  OAI222D0 U7963 ( .A1(n25003), .A2(n3606), .B1(n25004), .B2(n3510), .C1(
        n25005), .C2(n3558), .ZN(n25216) );
  OAI222D0 U7964 ( .A1(n24965), .A2(n2598), .B1(n25006), .B2(n3654), .C1(
        n25007), .C2(n3702), .ZN(n25215) );
  NR4D0 U7965 ( .A1(n25219), .A2(n25220), .A3(n25221), .A4(n25222), .ZN(n25203) );
  OAI22D0 U7966 ( .A1(n25012), .A2(n5142), .B1(n24966), .B2(n2310), .ZN(n25222) );
  OAI222D0 U7967 ( .A1(n24925), .A2(n3078), .B1(n24923), .B2(n2982), .C1(
        n24960), .C2(n2886), .ZN(n25221) );
  OAI222D0 U7968 ( .A1(n25013), .A2(n5526), .B1(n25014), .B2(n5574), .C1(
        n24924), .C2(n3030), .ZN(n25220) );
  OAI222D0 U7969 ( .A1(n25015), .A2(n6102), .B1(n25016), .B2(n6006), .C1(
        n25017), .C2(n6150), .ZN(n25219) );
  INR4D0 U7970 ( .A1(n25223), .B1(n25224), .B2(n25225), .B3(n25226), .ZN(
        n25201) );
  OAI222D0 U7971 ( .A1(n25022), .A2(n5478), .B1(n25023), .B2(n6342), .C1(
        n25024), .C2(n5430), .ZN(n25226) );
  OAI222D0 U7972 ( .A1(n25025), .A2(n4518), .B1(n25026), .B2(n24571), .C1(
        n25027), .C2(n5622), .ZN(n25225) );
  OR4D0 U7973 ( .A1(n25227), .A2(n25228), .A3(n25229), .A4(n25230), .Z(n25224)
         );
  OAI222D0 U7974 ( .A1(n25032), .A2(n4614), .B1(n25033), .B2(n5334), .C1(
        n25034), .C2(n6246), .ZN(n25230) );
  OAI222D0 U7975 ( .A1(n25035), .A2(n6198), .B1(n25036), .B2(n4566), .C1(
        n25037), .C2(n5382), .ZN(n25229) );
  OAI22D0 U7976 ( .A1(n27055), .A2(n25038), .B1(n27054), .B2(n25039), .ZN(
        n25228) );
  OAI222D0 U7977 ( .A1(n24906), .A2(n25040), .B1(n25041), .B2(n5862), .C1(
        n25042), .C2(n5814), .ZN(n25227) );
  CKND0 U7978 ( .I(\Mem[44][4] ), .ZN(n24906) );
  AOI221D0 U7979 ( .A1(n27052), .A2(n25043), .B1(n27053), .B2(n25044), .C(
        n25231), .ZN(n25223) );
  OAI222D0 U7980 ( .A1(n25046), .A2(n6054), .B1(n24907), .B2(n25047), .C1(
        n25048), .C2(n4710), .ZN(n25231) );
  CKND0 U7981 ( .I(\Mem[45][4] ), .ZN(n24907) );
  NR4D0 U7982 ( .A1(n25232), .A2(n25233), .A3(n25234), .A4(n25235), .ZN(n25200) );
  OAI22D0 U7983 ( .A1(n25053), .A2(n5910), .B1(n25054), .B2(n5718), .ZN(n25235) );
  OAI222D0 U7984 ( .A1(n25055), .A2(n3846), .B1(n25056), .B2(n3894), .C1(
        n25057), .C2(n5958), .ZN(n25234) );
  OAI222D0 U7985 ( .A1(n25058), .A2(n3990), .B1(n25059), .B2(n4038), .C1(
        n25060), .C2(n3942), .ZN(n25233) );
  OAI222D0 U7986 ( .A1(n25061), .A2(n4134), .B1(n25062), .B2(n4182), .C1(
        n25063), .C2(n4086), .ZN(n25232) );
  NR4D0 U7987 ( .A1(n25236), .A2(n25237), .A3(n25238), .A4(n25239), .ZN(n25199) );
  OAI22D0 U7988 ( .A1(n25068), .A2(n2406), .B1(n25069), .B2(n2934), .ZN(n25239) );
  OAI222D0 U7989 ( .A1(n25070), .A2(n2502), .B1(n25071), .B2(n4326), .C1(
        n25072), .C2(n2646), .ZN(n25238) );
  OAI222D0 U7990 ( .A1(n25073), .A2(n4278), .B1(n24930), .B2(n3318), .C1(
        n25074), .C2(n4230), .ZN(n25237) );
  OAI222D0 U7991 ( .A1(n24932), .A2(n3414), .B1(n25075), .B2(n4854), .C1(
        n24931), .C2(n3366), .ZN(n25236) );
  ND4D0 U7992 ( .A1(n25240), .A2(n25241), .A3(n25242), .A4(n25243), .ZN(n2213)
         );
  AN4D0 U7993 ( .A1(n25244), .A2(n25245), .A3(n25246), .A4(n25247), .Z(n25243)
         );
  NR4D0 U7994 ( .A1(n25248), .A2(n25249), .A3(n25250), .A4(n25251), .ZN(n25247) );
  OAI222D0 U7995 ( .A1(n24979), .A2(n15469), .B1(n24980), .B2(n4469), .C1(
        n24964), .C2(n2261), .ZN(n25251) );
  OAI222D0 U7996 ( .A1(n24920), .A2(n2549), .B1(n24981), .B2(n5189), .C1(
        n24963), .C2(n2453), .ZN(n25250) );
  OAI222D0 U7997 ( .A1(n24982), .A2(n4949), .B1(n24983), .B2(n4997), .C1(
        n24984), .C2(n4901), .ZN(n25249) );
  OAI222D0 U7998 ( .A1(n24985), .A2(n4421), .B1(n24986), .B2(n3797), .C1(
        n24987), .C2(n4373), .ZN(n25248) );
  NR4D0 U7999 ( .A1(n25252), .A2(n25253), .A3(n25254), .A4(n25255), .ZN(n25246) );
  OAI22D0 U8000 ( .A1(n24922), .A2(n2837), .B1(n24992), .B2(n3749), .ZN(n25255) );
  OAI222D0 U8001 ( .A1(n24993), .A2(n17941), .B1(n24962), .B2(n2789), .C1(
        n24994), .C2(n17942), .ZN(n25254) );
  OAI222D0 U8002 ( .A1(n24995), .A2(n5237), .B1(n24961), .B2(n2693), .C1(
        n24921), .C2(n2741), .ZN(n25253) );
  OAI222D0 U8003 ( .A1(n24927), .A2(n3173), .B1(n24996), .B2(n4805), .C1(
        n24997), .C2(n15468), .ZN(n25252) );
  NR4D0 U8004 ( .A1(n25256), .A2(n25257), .A3(n25258), .A4(n25259), .ZN(n25245) );
  OAI22D0 U8005 ( .A1(n24928), .A2(n3221), .B1(n24926), .B2(n3125), .ZN(n25259) );
  OAI222D0 U8006 ( .A1(n25002), .A2(n3461), .B1(n24929), .B2(n3269), .C1(
        n24933), .C2(n2357), .ZN(n25258) );
  OAI222D0 U8007 ( .A1(n25003), .A2(n3605), .B1(n25004), .B2(n3509), .C1(
        n25005), .C2(n3557), .ZN(n25257) );
  OAI222D0 U8008 ( .A1(n24965), .A2(n2597), .B1(n25006), .B2(n3653), .C1(
        n25007), .C2(n3701), .ZN(n25256) );
  NR4D0 U8009 ( .A1(n25260), .A2(n25261), .A3(n25262), .A4(n25263), .ZN(n25244) );
  OAI22D0 U8010 ( .A1(n25012), .A2(n5141), .B1(n24966), .B2(n2309), .ZN(n25263) );
  OAI222D0 U8011 ( .A1(n24925), .A2(n3077), .B1(n24923), .B2(n2981), .C1(
        n24960), .C2(n2885), .ZN(n25262) );
  OAI222D0 U8012 ( .A1(n25013), .A2(n5525), .B1(n25014), .B2(n5573), .C1(
        n24924), .C2(n3029), .ZN(n25261) );
  OAI222D0 U8013 ( .A1(n25015), .A2(n6101), .B1(n25016), .B2(n6005), .C1(
        n25017), .C2(n6149), .ZN(n25260) );
  INR4D0 U8014 ( .A1(n25264), .B1(n25265), .B2(n25266), .B3(n25267), .ZN(
        n25242) );
  OAI222D0 U8015 ( .A1(n25022), .A2(n5477), .B1(n25023), .B2(n6341), .C1(
        n25024), .C2(n5429), .ZN(n25267) );
  OAI222D0 U8016 ( .A1(n25025), .A2(n4517), .B1(n25026), .B2(n24574), .C1(
        n25027), .C2(n5621), .ZN(n25266) );
  OR4D0 U8017 ( .A1(n25268), .A2(n25269), .A3(n25270), .A4(n25271), .Z(n25265)
         );
  OAI222D0 U8018 ( .A1(n25032), .A2(n4613), .B1(n25033), .B2(n5333), .C1(
        n25034), .C2(n6245), .ZN(n25271) );
  OAI222D0 U8019 ( .A1(n25035), .A2(n6197), .B1(n25036), .B2(n4565), .C1(
        n25037), .C2(n5381), .ZN(n25270) );
  OAI22D0 U8020 ( .A1(n27059), .A2(n25038), .B1(n27058), .B2(n25039), .ZN(
        n25269) );
  OAI222D0 U8021 ( .A1(n24904), .A2(n25040), .B1(n25041), .B2(n5861), .C1(
        n25042), .C2(n5813), .ZN(n25268) );
  CKND0 U8022 ( .I(\Mem[44][5] ), .ZN(n24904) );
  AOI221D0 U8023 ( .A1(n27056), .A2(n25043), .B1(n27057), .B2(n25044), .C(
        n25272), .ZN(n25264) );
  OAI222D0 U8024 ( .A1(n25046), .A2(n6053), .B1(n24905), .B2(n25047), .C1(
        n25048), .C2(n4709), .ZN(n25272) );
  CKND0 U8025 ( .I(\Mem[45][5] ), .ZN(n24905) );
  NR4D0 U8026 ( .A1(n25273), .A2(n25274), .A3(n25275), .A4(n25276), .ZN(n25241) );
  OAI22D0 U8027 ( .A1(n25053), .A2(n5909), .B1(n25054), .B2(n5717), .ZN(n25276) );
  OAI222D0 U8028 ( .A1(n25055), .A2(n3845), .B1(n25056), .B2(n3893), .C1(
        n25057), .C2(n5957), .ZN(n25275) );
  OAI222D0 U8029 ( .A1(n25058), .A2(n3989), .B1(n25059), .B2(n4037), .C1(
        n25060), .C2(n3941), .ZN(n25274) );
  OAI222D0 U8030 ( .A1(n25061), .A2(n4133), .B1(n25062), .B2(n4181), .C1(
        n25063), .C2(n4085), .ZN(n25273) );
  NR4D0 U8031 ( .A1(n25277), .A2(n25278), .A3(n25279), .A4(n25280), .ZN(n25240) );
  OAI22D0 U8032 ( .A1(n25068), .A2(n2405), .B1(n25069), .B2(n2933), .ZN(n25280) );
  OAI222D0 U8033 ( .A1(n25070), .A2(n2501), .B1(n25071), .B2(n4325), .C1(
        n25072), .C2(n2645), .ZN(n25279) );
  OAI222D0 U8034 ( .A1(n25073), .A2(n4277), .B1(n24930), .B2(n3317), .C1(
        n25074), .C2(n4229), .ZN(n25278) );
  OAI222D0 U8035 ( .A1(n24932), .A2(n3413), .B1(n25075), .B2(n4853), .C1(
        n24931), .C2(n3365), .ZN(n25277) );
  ND4D0 U8036 ( .A1(n25281), .A2(n25282), .A3(n25283), .A4(n25284), .ZN(n2212)
         );
  AN4D0 U8037 ( .A1(n25285), .A2(n25286), .A3(n25287), .A4(n25288), .Z(n25284)
         );
  NR4D0 U8038 ( .A1(n25289), .A2(n25290), .A3(n25291), .A4(n25292), .ZN(n25288) );
  OAI222D0 U8039 ( .A1(n24979), .A2(n15473), .B1(n24980), .B2(n4468), .C1(
        n24964), .C2(n2260), .ZN(n25292) );
  OAI222D0 U8040 ( .A1(n24920), .A2(n2548), .B1(n24981), .B2(n5188), .C1(
        n24963), .C2(n2452), .ZN(n25291) );
  OAI222D0 U8041 ( .A1(n24982), .A2(n4948), .B1(n24983), .B2(n4996), .C1(
        n24984), .C2(n4900), .ZN(n25290) );
  OAI222D0 U8042 ( .A1(n24985), .A2(n4420), .B1(n24986), .B2(n3796), .C1(
        n24987), .C2(n4372), .ZN(n25289) );
  NR4D0 U8043 ( .A1(n25293), .A2(n25294), .A3(n25295), .A4(n25296), .ZN(n25287) );
  OAI22D0 U8044 ( .A1(n24922), .A2(n2836), .B1(n24992), .B2(n3748), .ZN(n25296) );
  OAI222D0 U8045 ( .A1(n24993), .A2(n17944), .B1(n24962), .B2(n2788), .C1(
        n24994), .C2(n17945), .ZN(n25295) );
  OAI222D0 U8046 ( .A1(n24995), .A2(n5236), .B1(n24961), .B2(n2692), .C1(
        n24921), .C2(n2740), .ZN(n25294) );
  OAI222D0 U8047 ( .A1(n24927), .A2(n3172), .B1(n24996), .B2(n4804), .C1(
        n24997), .C2(n15472), .ZN(n25293) );
  NR4D0 U8048 ( .A1(n25297), .A2(n25298), .A3(n25299), .A4(n25300), .ZN(n25286) );
  OAI22D0 U8049 ( .A1(n24928), .A2(n3220), .B1(n24926), .B2(n3124), .ZN(n25300) );
  OAI222D0 U8050 ( .A1(n25002), .A2(n3460), .B1(n24929), .B2(n3268), .C1(
        n24933), .C2(n2356), .ZN(n25299) );
  OAI222D0 U8051 ( .A1(n25003), .A2(n3604), .B1(n25004), .B2(n3508), .C1(
        n25005), .C2(n3556), .ZN(n25298) );
  OAI222D0 U8052 ( .A1(n24965), .A2(n2596), .B1(n25006), .B2(n3652), .C1(
        n25007), .C2(n3700), .ZN(n25297) );
  NR4D0 U8053 ( .A1(n25301), .A2(n25302), .A3(n25303), .A4(n25304), .ZN(n25285) );
  OAI22D0 U8054 ( .A1(n25012), .A2(n5140), .B1(n24966), .B2(n2308), .ZN(n25304) );
  OAI222D0 U8055 ( .A1(n24925), .A2(n3076), .B1(n24923), .B2(n2980), .C1(
        n24960), .C2(n2884), .ZN(n25303) );
  OAI222D0 U8056 ( .A1(n25013), .A2(n5524), .B1(n25014), .B2(n5572), .C1(
        n24924), .C2(n3028), .ZN(n25302) );
  OAI222D0 U8057 ( .A1(n25015), .A2(n6100), .B1(n25016), .B2(n6004), .C1(
        n25017), .C2(n6148), .ZN(n25301) );
  INR4D0 U8058 ( .A1(n25305), .B1(n25306), .B2(n25307), .B3(n25308), .ZN(
        n25283) );
  OAI222D0 U8059 ( .A1(n25022), .A2(n5476), .B1(n25023), .B2(n6340), .C1(
        n25024), .C2(n5428), .ZN(n25308) );
  OAI222D0 U8060 ( .A1(n25025), .A2(n4516), .B1(n25026), .B2(n24577), .C1(
        n25027), .C2(n5620), .ZN(n25307) );
  OR4D0 U8061 ( .A1(n25309), .A2(n25310), .A3(n25311), .A4(n25312), .Z(n25306)
         );
  OAI222D0 U8062 ( .A1(n25032), .A2(n4612), .B1(n25033), .B2(n5332), .C1(
        n25034), .C2(n6244), .ZN(n25312) );
  OAI222D0 U8063 ( .A1(n25035), .A2(n6196), .B1(n25036), .B2(n4564), .C1(
        n25037), .C2(n5380), .ZN(n25311) );
  OAI22D0 U8064 ( .A1(n27063), .A2(n25038), .B1(n27062), .B2(n25039), .ZN(
        n25310) );
  OAI222D0 U8065 ( .A1(n24902), .A2(n25040), .B1(n25041), .B2(n5860), .C1(
        n25042), .C2(n5812), .ZN(n25309) );
  CKND0 U8066 ( .I(\Mem[44][6] ), .ZN(n24902) );
  AOI221D0 U8067 ( .A1(n27060), .A2(n25043), .B1(n27061), .B2(n25044), .C(
        n25313), .ZN(n25305) );
  OAI222D0 U8068 ( .A1(n25046), .A2(n6052), .B1(n24903), .B2(n25047), .C1(
        n25048), .C2(n4708), .ZN(n25313) );
  CKND0 U8069 ( .I(\Mem[45][6] ), .ZN(n24903) );
  NR4D0 U8070 ( .A1(n25314), .A2(n25315), .A3(n25316), .A4(n25317), .ZN(n25282) );
  OAI22D0 U8071 ( .A1(n25053), .A2(n5908), .B1(n25054), .B2(n5716), .ZN(n25317) );
  OAI222D0 U8072 ( .A1(n25055), .A2(n3844), .B1(n25056), .B2(n3892), .C1(
        n25057), .C2(n5956), .ZN(n25316) );
  OAI222D0 U8073 ( .A1(n25058), .A2(n3988), .B1(n25059), .B2(n4036), .C1(
        n25060), .C2(n3940), .ZN(n25315) );
  OAI222D0 U8074 ( .A1(n25061), .A2(n4132), .B1(n25062), .B2(n4180), .C1(
        n25063), .C2(n4084), .ZN(n25314) );
  NR4D0 U8075 ( .A1(n25318), .A2(n25319), .A3(n25320), .A4(n25321), .ZN(n25281) );
  OAI22D0 U8076 ( .A1(n25068), .A2(n2404), .B1(n25069), .B2(n2932), .ZN(n25321) );
  OAI222D0 U8077 ( .A1(n25070), .A2(n2500), .B1(n25071), .B2(n4324), .C1(
        n25072), .C2(n2644), .ZN(n25320) );
  OAI222D0 U8078 ( .A1(n25073), .A2(n4276), .B1(n24930), .B2(n3316), .C1(
        n25074), .C2(n4228), .ZN(n25319) );
  OAI222D0 U8079 ( .A1(n24932), .A2(n3412), .B1(n25075), .B2(n4852), .C1(
        n24931), .C2(n3364), .ZN(n25318) );
  ND4D0 U8080 ( .A1(n25322), .A2(n25323), .A3(n25324), .A4(n25325), .ZN(n2211)
         );
  AN4D0 U8081 ( .A1(n25326), .A2(n25327), .A3(n25328), .A4(n25329), .Z(n25325)
         );
  NR4D0 U8082 ( .A1(n25330), .A2(n25331), .A3(n25332), .A4(n25333), .ZN(n25329) );
  OAI222D0 U8083 ( .A1(n24979), .A2(n15477), .B1(n24980), .B2(n4467), .C1(
        n24964), .C2(n2259), .ZN(n25333) );
  OAI222D0 U8084 ( .A1(n24920), .A2(n2547), .B1(n24981), .B2(n5187), .C1(
        n24963), .C2(n2451), .ZN(n25332) );
  OAI222D0 U8085 ( .A1(n24982), .A2(n4947), .B1(n24983), .B2(n4995), .C1(
        n24984), .C2(n4899), .ZN(n25331) );
  OAI222D0 U8086 ( .A1(n24985), .A2(n4419), .B1(n24986), .B2(n3795), .C1(
        n24987), .C2(n4371), .ZN(n25330) );
  NR4D0 U8087 ( .A1(n25334), .A2(n25335), .A3(n25336), .A4(n25337), .ZN(n25328) );
  OAI22D0 U8088 ( .A1(n24922), .A2(n2835), .B1(n24992), .B2(n3747), .ZN(n25337) );
  OAI222D0 U8089 ( .A1(n24993), .A2(n17947), .B1(n24962), .B2(n2787), .C1(
        n24994), .C2(n17948), .ZN(n25336) );
  OAI222D0 U8090 ( .A1(n24995), .A2(n5235), .B1(n24961), .B2(n2691), .C1(
        n24921), .C2(n2739), .ZN(n25335) );
  OAI222D0 U8091 ( .A1(n24927), .A2(n3171), .B1(n24996), .B2(n4803), .C1(
        n24997), .C2(n15476), .ZN(n25334) );
  NR4D0 U8092 ( .A1(n25338), .A2(n25339), .A3(n25340), .A4(n25341), .ZN(n25327) );
  OAI22D0 U8093 ( .A1(n24928), .A2(n3219), .B1(n24926), .B2(n3123), .ZN(n25341) );
  OAI222D0 U8094 ( .A1(n25002), .A2(n3459), .B1(n24929), .B2(n3267), .C1(
        n24933), .C2(n2355), .ZN(n25340) );
  OAI222D0 U8095 ( .A1(n25003), .A2(n3603), .B1(n25004), .B2(n3507), .C1(
        n25005), .C2(n3555), .ZN(n25339) );
  OAI222D0 U8096 ( .A1(n24965), .A2(n2595), .B1(n25006), .B2(n3651), .C1(
        n25007), .C2(n3699), .ZN(n25338) );
  NR4D0 U8097 ( .A1(n25342), .A2(n25343), .A3(n25344), .A4(n25345), .ZN(n25326) );
  OAI22D0 U8098 ( .A1(n25012), .A2(n5139), .B1(n24966), .B2(n2307), .ZN(n25345) );
  OAI222D0 U8099 ( .A1(n24925), .A2(n3075), .B1(n24923), .B2(n2979), .C1(
        n24960), .C2(n2883), .ZN(n25344) );
  OAI222D0 U8100 ( .A1(n25013), .A2(n5523), .B1(n25014), .B2(n5571), .C1(
        n24924), .C2(n3027), .ZN(n25343) );
  OAI222D0 U8101 ( .A1(n25015), .A2(n6099), .B1(n25016), .B2(n6003), .C1(
        n25017), .C2(n6147), .ZN(n25342) );
  INR4D0 U8102 ( .A1(n25346), .B1(n25347), .B2(n25348), .B3(n25349), .ZN(
        n25324) );
  OAI222D0 U8103 ( .A1(n25022), .A2(n5475), .B1(n25023), .B2(n6339), .C1(
        n25024), .C2(n5427), .ZN(n25349) );
  OAI222D0 U8104 ( .A1(n25025), .A2(n4515), .B1(n25026), .B2(n24580), .C1(
        n25027), .C2(n5619), .ZN(n25348) );
  OR4D0 U8105 ( .A1(n25350), .A2(n25351), .A3(n25352), .A4(n25353), .Z(n25347)
         );
  OAI222D0 U8106 ( .A1(n25032), .A2(n4611), .B1(n25033), .B2(n5331), .C1(
        n25034), .C2(n6243), .ZN(n25353) );
  OAI222D0 U8107 ( .A1(n25035), .A2(n6195), .B1(n25036), .B2(n4563), .C1(
        n25037), .C2(n5379), .ZN(n25352) );
  OAI22D0 U8108 ( .A1(n27067), .A2(n25038), .B1(n27066), .B2(n25039), .ZN(
        n25351) );
  OAI222D0 U8109 ( .A1(n24900), .A2(n25040), .B1(n25041), .B2(n5859), .C1(
        n25042), .C2(n5811), .ZN(n25350) );
  CKND0 U8110 ( .I(\Mem[44][7] ), .ZN(n24900) );
  AOI221D0 U8111 ( .A1(n27064), .A2(n25043), .B1(n27065), .B2(n25044), .C(
        n25354), .ZN(n25346) );
  OAI222D0 U8112 ( .A1(n25046), .A2(n6051), .B1(n24901), .B2(n25047), .C1(
        n25048), .C2(n4707), .ZN(n25354) );
  CKND0 U8113 ( .I(\Mem[45][7] ), .ZN(n24901) );
  NR4D0 U8114 ( .A1(n25355), .A2(n25356), .A3(n25357), .A4(n25358), .ZN(n25323) );
  OAI22D0 U8115 ( .A1(n25053), .A2(n5907), .B1(n25054), .B2(n5715), .ZN(n25358) );
  OAI222D0 U8116 ( .A1(n25055), .A2(n3843), .B1(n25056), .B2(n3891), .C1(
        n25057), .C2(n5955), .ZN(n25357) );
  OAI222D0 U8117 ( .A1(n25058), .A2(n3987), .B1(n25059), .B2(n4035), .C1(
        n25060), .C2(n3939), .ZN(n25356) );
  OAI222D0 U8118 ( .A1(n25061), .A2(n4131), .B1(n25062), .B2(n4179), .C1(
        n25063), .C2(n4083), .ZN(n25355) );
  NR4D0 U8119 ( .A1(n25359), .A2(n25360), .A3(n25361), .A4(n25362), .ZN(n25322) );
  OAI22D0 U8120 ( .A1(n25068), .A2(n2403), .B1(n25069), .B2(n2931), .ZN(n25362) );
  OAI222D0 U8121 ( .A1(n25070), .A2(n2499), .B1(n25071), .B2(n4323), .C1(
        n25072), .C2(n2643), .ZN(n25361) );
  OAI222D0 U8122 ( .A1(n25073), .A2(n4275), .B1(n24930), .B2(n3315), .C1(
        n25074), .C2(n4227), .ZN(n25360) );
  OAI222D0 U8123 ( .A1(n24932), .A2(n3411), .B1(n25075), .B2(n4851), .C1(
        n24931), .C2(n3363), .ZN(n25359) );
  ND4D0 U8124 ( .A1(n25363), .A2(n25364), .A3(n25365), .A4(n25366), .ZN(n2210)
         );
  AN4D0 U8125 ( .A1(n25367), .A2(n25368), .A3(n25369), .A4(n25370), .Z(n25366)
         );
  NR4D0 U8126 ( .A1(n25371), .A2(n25372), .A3(n25373), .A4(n25374), .ZN(n25370) );
  OAI222D0 U8127 ( .A1(n24979), .A2(n15481), .B1(n24980), .B2(n4466), .C1(
        n24964), .C2(n2258), .ZN(n25374) );
  OAI222D0 U8128 ( .A1(n24920), .A2(n2546), .B1(n24981), .B2(n5186), .C1(
        n24963), .C2(n2450), .ZN(n25373) );
  OAI222D0 U8129 ( .A1(n24982), .A2(n4946), .B1(n24983), .B2(n4994), .C1(
        n24984), .C2(n4898), .ZN(n25372) );
  OAI222D0 U8130 ( .A1(n24985), .A2(n4418), .B1(n24986), .B2(n3794), .C1(
        n24987), .C2(n4370), .ZN(n25371) );
  NR4D0 U8131 ( .A1(n25375), .A2(n25376), .A3(n25377), .A4(n25378), .ZN(n25369) );
  OAI22D0 U8132 ( .A1(n24922), .A2(n2834), .B1(n24992), .B2(n3746), .ZN(n25378) );
  OAI222D0 U8133 ( .A1(n24993), .A2(n17950), .B1(n24962), .B2(n2786), .C1(
        n24994), .C2(n17951), .ZN(n25377) );
  OAI222D0 U8134 ( .A1(n24995), .A2(n5234), .B1(n24961), .B2(n2690), .C1(
        n24921), .C2(n2738), .ZN(n25376) );
  OAI222D0 U8135 ( .A1(n24927), .A2(n3170), .B1(n24996), .B2(n4802), .C1(
        n24997), .C2(n15480), .ZN(n25375) );
  NR4D0 U8136 ( .A1(n25379), .A2(n25380), .A3(n25381), .A4(n25382), .ZN(n25368) );
  OAI22D0 U8137 ( .A1(n24928), .A2(n3218), .B1(n24926), .B2(n3122), .ZN(n25382) );
  OAI222D0 U8138 ( .A1(n25002), .A2(n3458), .B1(n24929), .B2(n3266), .C1(
        n24933), .C2(n2354), .ZN(n25381) );
  OAI222D0 U8139 ( .A1(n25003), .A2(n3602), .B1(n25004), .B2(n3506), .C1(
        n25005), .C2(n3554), .ZN(n25380) );
  OAI222D0 U8140 ( .A1(n24965), .A2(n2594), .B1(n25006), .B2(n3650), .C1(
        n25007), .C2(n3698), .ZN(n25379) );
  NR4D0 U8141 ( .A1(n25383), .A2(n25384), .A3(n25385), .A4(n25386), .ZN(n25367) );
  OAI22D0 U8142 ( .A1(n25012), .A2(n5138), .B1(n24966), .B2(n2306), .ZN(n25386) );
  OAI222D0 U8143 ( .A1(n24925), .A2(n3074), .B1(n24923), .B2(n2978), .C1(
        n24960), .C2(n2882), .ZN(n25385) );
  OAI222D0 U8144 ( .A1(n25013), .A2(n5522), .B1(n25014), .B2(n5570), .C1(
        n24924), .C2(n3026), .ZN(n25384) );
  OAI222D0 U8145 ( .A1(n25015), .A2(n6098), .B1(n25016), .B2(n6002), .C1(
        n25017), .C2(n6146), .ZN(n25383) );
  INR4D0 U8146 ( .A1(n25387), .B1(n25388), .B2(n25389), .B3(n25390), .ZN(
        n25365) );
  OAI222D0 U8147 ( .A1(n25022), .A2(n5474), .B1(n25023), .B2(n6338), .C1(
        n25024), .C2(n5426), .ZN(n25390) );
  OAI222D0 U8148 ( .A1(n25025), .A2(n4514), .B1(n25026), .B2(n24583), .C1(
        n25027), .C2(n5618), .ZN(n25389) );
  OR4D0 U8149 ( .A1(n25391), .A2(n25392), .A3(n25393), .A4(n25394), .Z(n25388)
         );
  OAI222D0 U8150 ( .A1(n25032), .A2(n4610), .B1(n25033), .B2(n5330), .C1(
        n25034), .C2(n6242), .ZN(n25394) );
  OAI222D0 U8151 ( .A1(n25035), .A2(n6194), .B1(n25036), .B2(n4562), .C1(
        n25037), .C2(n5378), .ZN(n25393) );
  OAI22D0 U8152 ( .A1(n27071), .A2(n25038), .B1(n27070), .B2(n25039), .ZN(
        n25392) );
  OAI222D0 U8153 ( .A1(n24898), .A2(n25040), .B1(n25041), .B2(n5858), .C1(
        n25042), .C2(n5810), .ZN(n25391) );
  CKND0 U8154 ( .I(\Mem[44][8] ), .ZN(n24898) );
  AOI221D0 U8155 ( .A1(n27068), .A2(n25043), .B1(n27069), .B2(n25044), .C(
        n25395), .ZN(n25387) );
  OAI222D0 U8156 ( .A1(n25046), .A2(n6050), .B1(n24899), .B2(n25047), .C1(
        n25048), .C2(n4706), .ZN(n25395) );
  CKND0 U8157 ( .I(\Mem[45][8] ), .ZN(n24899) );
  NR4D0 U8158 ( .A1(n25396), .A2(n25397), .A3(n25398), .A4(n25399), .ZN(n25364) );
  OAI22D0 U8159 ( .A1(n25053), .A2(n5906), .B1(n25054), .B2(n5714), .ZN(n25399) );
  OAI222D0 U8160 ( .A1(n25055), .A2(n3842), .B1(n25056), .B2(n3890), .C1(
        n25057), .C2(n5954), .ZN(n25398) );
  OAI222D0 U8161 ( .A1(n25058), .A2(n3986), .B1(n25059), .B2(n4034), .C1(
        n25060), .C2(n3938), .ZN(n25397) );
  OAI222D0 U8162 ( .A1(n25061), .A2(n4130), .B1(n25062), .B2(n4178), .C1(
        n25063), .C2(n4082), .ZN(n25396) );
  NR4D0 U8163 ( .A1(n25400), .A2(n25401), .A3(n25402), .A4(n25403), .ZN(n25363) );
  OAI22D0 U8164 ( .A1(n25068), .A2(n2402), .B1(n25069), .B2(n2930), .ZN(n25403) );
  OAI222D0 U8165 ( .A1(n25070), .A2(n2498), .B1(n25071), .B2(n4322), .C1(
        n25072), .C2(n2642), .ZN(n25402) );
  OAI222D0 U8166 ( .A1(n25073), .A2(n4274), .B1(n24930), .B2(n3314), .C1(
        n25074), .C2(n4226), .ZN(n25401) );
  OAI222D0 U8167 ( .A1(n24932), .A2(n3410), .B1(n25075), .B2(n4850), .C1(
        n24931), .C2(n3362), .ZN(n25400) );
  ND4D0 U8168 ( .A1(n25404), .A2(n25405), .A3(n25406), .A4(n25407), .ZN(n2208)
         );
  AN4D0 U8169 ( .A1(n25408), .A2(n25409), .A3(n25410), .A4(n25411), .Z(n25407)
         );
  NR4D0 U8170 ( .A1(n25412), .A2(n25413), .A3(n25414), .A4(n25415), .ZN(n25411) );
  OAI222D0 U8171 ( .A1(n24979), .A2(n15485), .B1(n24980), .B2(n4465), .C1(
        n24964), .C2(n2257), .ZN(n25415) );
  OAI222D0 U8172 ( .A1(n24920), .A2(n2545), .B1(n24981), .B2(n5185), .C1(
        n24963), .C2(n2449), .ZN(n25414) );
  OAI222D0 U8173 ( .A1(n24982), .A2(n4945), .B1(n24983), .B2(n4993), .C1(
        n24984), .C2(n4897), .ZN(n25413) );
  OAI222D0 U8174 ( .A1(n24985), .A2(n4417), .B1(n24986), .B2(n3793), .C1(
        n24987), .C2(n4369), .ZN(n25412) );
  NR4D0 U8175 ( .A1(n25416), .A2(n25417), .A3(n25418), .A4(n25419), .ZN(n25410) );
  OAI22D0 U8176 ( .A1(n24922), .A2(n2833), .B1(n24992), .B2(n3745), .ZN(n25419) );
  OAI222D0 U8177 ( .A1(n24993), .A2(n17953), .B1(n24962), .B2(n2785), .C1(
        n24994), .C2(n17954), .ZN(n25418) );
  OAI222D0 U8178 ( .A1(n24995), .A2(n5233), .B1(n24961), .B2(n2689), .C1(
        n24921), .C2(n2737), .ZN(n25417) );
  OAI222D0 U8179 ( .A1(n24927), .A2(n3169), .B1(n24996), .B2(n4801), .C1(
        n24997), .C2(n15484), .ZN(n25416) );
  NR4D0 U8180 ( .A1(n25420), .A2(n25421), .A3(n25422), .A4(n25423), .ZN(n25409) );
  OAI22D0 U8181 ( .A1(n24928), .A2(n3217), .B1(n24926), .B2(n3121), .ZN(n25423) );
  OAI222D0 U8182 ( .A1(n25002), .A2(n3457), .B1(n24929), .B2(n3265), .C1(
        n24933), .C2(n2353), .ZN(n25422) );
  OAI222D0 U8183 ( .A1(n25003), .A2(n3601), .B1(n25004), .B2(n3505), .C1(
        n25005), .C2(n3553), .ZN(n25421) );
  OAI222D0 U8184 ( .A1(n24965), .A2(n2593), .B1(n25006), .B2(n3649), .C1(
        n25007), .C2(n3697), .ZN(n25420) );
  NR4D0 U8185 ( .A1(n25424), .A2(n25425), .A3(n25426), .A4(n25427), .ZN(n25408) );
  OAI22D0 U8186 ( .A1(n25012), .A2(n5137), .B1(n24966), .B2(n2305), .ZN(n25427) );
  OAI222D0 U8187 ( .A1(n24925), .A2(n3073), .B1(n24923), .B2(n2977), .C1(
        n24960), .C2(n2881), .ZN(n25426) );
  OAI222D0 U8188 ( .A1(n25013), .A2(n5521), .B1(n25014), .B2(n5569), .C1(
        n24924), .C2(n3025), .ZN(n25425) );
  OAI222D0 U8189 ( .A1(n25015), .A2(n6097), .B1(n25016), .B2(n6001), .C1(
        n25017), .C2(n6145), .ZN(n25424) );
  INR4D0 U8190 ( .A1(n25428), .B1(n25429), .B2(n25430), .B3(n25431), .ZN(
        n25406) );
  OAI222D0 U8191 ( .A1(n25022), .A2(n5473), .B1(n25023), .B2(n6337), .C1(
        n25024), .C2(n5425), .ZN(n25431) );
  OAI222D0 U8192 ( .A1(n25025), .A2(n4513), .B1(n25026), .B2(n24586), .C1(
        n25027), .C2(n5617), .ZN(n25430) );
  OR4D0 U8193 ( .A1(n25432), .A2(n25433), .A3(n25434), .A4(n25435), .Z(n25429)
         );
  OAI222D0 U8194 ( .A1(n25032), .A2(n4609), .B1(n25033), .B2(n5329), .C1(
        n25034), .C2(n6241), .ZN(n25435) );
  OAI222D0 U8195 ( .A1(n25035), .A2(n6193), .B1(n25036), .B2(n4561), .C1(
        n25037), .C2(n5377), .ZN(n25434) );
  OAI22D0 U8196 ( .A1(n27075), .A2(n25038), .B1(n27074), .B2(n25039), .ZN(
        n25433) );
  OAI222D0 U8197 ( .A1(n24896), .A2(n25040), .B1(n25041), .B2(n5857), .C1(
        n25042), .C2(n5809), .ZN(n25432) );
  CKND0 U8198 ( .I(\Mem[44][9] ), .ZN(n24896) );
  AOI221D0 U8199 ( .A1(n27072), .A2(n25043), .B1(n27073), .B2(n25044), .C(
        n25436), .ZN(n25428) );
  OAI222D0 U8200 ( .A1(n25046), .A2(n6049), .B1(n24897), .B2(n25047), .C1(
        n25048), .C2(n4705), .ZN(n25436) );
  CKND0 U8201 ( .I(\Mem[45][9] ), .ZN(n24897) );
  NR4D0 U8202 ( .A1(n25437), .A2(n25438), .A3(n25439), .A4(n25440), .ZN(n25405) );
  OAI22D0 U8203 ( .A1(n25053), .A2(n5905), .B1(n25054), .B2(n5713), .ZN(n25440) );
  OAI222D0 U8204 ( .A1(n25055), .A2(n3841), .B1(n25056), .B2(n3889), .C1(
        n25057), .C2(n5953), .ZN(n25439) );
  OAI222D0 U8205 ( .A1(n25058), .A2(n3985), .B1(n25059), .B2(n4033), .C1(
        n25060), .C2(n3937), .ZN(n25438) );
  OAI222D0 U8206 ( .A1(n25061), .A2(n4129), .B1(n25062), .B2(n4177), .C1(
        n25063), .C2(n4081), .ZN(n25437) );
  NR4D0 U8207 ( .A1(n25441), .A2(n25442), .A3(n25443), .A4(n25444), .ZN(n25404) );
  OAI22D0 U8208 ( .A1(n25068), .A2(n2401), .B1(n25069), .B2(n2929), .ZN(n25444) );
  OAI222D0 U8209 ( .A1(n25070), .A2(n2497), .B1(n25071), .B2(n4321), .C1(
        n25072), .C2(n2641), .ZN(n25443) );
  OAI222D0 U8210 ( .A1(n25073), .A2(n4273), .B1(n24930), .B2(n3313), .C1(
        n25074), .C2(n4225), .ZN(n25442) );
  OAI222D0 U8211 ( .A1(n24932), .A2(n3409), .B1(n25075), .B2(n4849), .C1(
        n24931), .C2(n3361), .ZN(n25441) );
  ND4D0 U8212 ( .A1(n25445), .A2(n25446), .A3(n25447), .A4(n25448), .ZN(n2207)
         );
  AN4D0 U8213 ( .A1(n25449), .A2(n25450), .A3(n25451), .A4(n25452), .Z(n25448)
         );
  NR4D0 U8214 ( .A1(n25453), .A2(n25454), .A3(n25455), .A4(n25456), .ZN(n25452) );
  OAI222D0 U8215 ( .A1(n24979), .A2(n15489), .B1(n24980), .B2(n4464), .C1(
        n24964), .C2(n2256), .ZN(n25456) );
  OAI222D0 U8216 ( .A1(n24920), .A2(n2544), .B1(n24981), .B2(n5184), .C1(
        n24963), .C2(n2448), .ZN(n25455) );
  OAI222D0 U8217 ( .A1(n24982), .A2(n4944), .B1(n24983), .B2(n4992), .C1(
        n24984), .C2(n4896), .ZN(n25454) );
  OAI222D0 U8218 ( .A1(n24985), .A2(n4416), .B1(n24986), .B2(n3792), .C1(
        n24987), .C2(n4368), .ZN(n25453) );
  NR4D0 U8219 ( .A1(n25457), .A2(n25458), .A3(n25459), .A4(n25460), .ZN(n25451) );
  OAI22D0 U8220 ( .A1(n24922), .A2(n2832), .B1(n24992), .B2(n3744), .ZN(n25460) );
  OAI222D0 U8221 ( .A1(n24993), .A2(n17956), .B1(n24962), .B2(n2784), .C1(
        n24994), .C2(n17957), .ZN(n25459) );
  OAI222D0 U8222 ( .A1(n24995), .A2(n5232), .B1(n24961), .B2(n2688), .C1(
        n24921), .C2(n2736), .ZN(n25458) );
  OAI222D0 U8223 ( .A1(n24927), .A2(n3168), .B1(n24996), .B2(n4800), .C1(
        n24997), .C2(n15488), .ZN(n25457) );
  NR4D0 U8224 ( .A1(n25461), .A2(n25462), .A3(n25463), .A4(n25464), .ZN(n25450) );
  OAI22D0 U8225 ( .A1(n24928), .A2(n3216), .B1(n24926), .B2(n3120), .ZN(n25464) );
  OAI222D0 U8226 ( .A1(n25002), .A2(n3456), .B1(n24929), .B2(n3264), .C1(
        n24933), .C2(n2352), .ZN(n25463) );
  OAI222D0 U8227 ( .A1(n25003), .A2(n3600), .B1(n25004), .B2(n3504), .C1(
        n25005), .C2(n3552), .ZN(n25462) );
  OAI222D0 U8228 ( .A1(n24965), .A2(n2592), .B1(n25006), .B2(n3648), .C1(
        n25007), .C2(n3696), .ZN(n25461) );
  NR4D0 U8229 ( .A1(n25465), .A2(n25466), .A3(n25467), .A4(n25468), .ZN(n25449) );
  OAI22D0 U8230 ( .A1(n25012), .A2(n5136), .B1(n24966), .B2(n2304), .ZN(n25468) );
  OAI222D0 U8231 ( .A1(n24925), .A2(n3072), .B1(n24923), .B2(n2976), .C1(
        n24960), .C2(n2880), .ZN(n25467) );
  OAI222D0 U8232 ( .A1(n25013), .A2(n5520), .B1(n25014), .B2(n5568), .C1(
        n24924), .C2(n3024), .ZN(n25466) );
  OAI222D0 U8233 ( .A1(n25015), .A2(n6096), .B1(n25016), .B2(n6000), .C1(
        n25017), .C2(n6144), .ZN(n25465) );
  INR4D0 U8234 ( .A1(n25469), .B1(n25470), .B2(n25471), .B3(n25472), .ZN(
        n25447) );
  OAI222D0 U8235 ( .A1(n25022), .A2(n5472), .B1(n25023), .B2(n6336), .C1(
        n25024), .C2(n5424), .ZN(n25472) );
  OAI222D0 U8236 ( .A1(n25025), .A2(n4512), .B1(n25026), .B2(n24589), .C1(
        n25027), .C2(n5616), .ZN(n25471) );
  OR4D0 U8237 ( .A1(n25473), .A2(n25474), .A3(n25475), .A4(n25476), .Z(n25470)
         );
  OAI222D0 U8238 ( .A1(n25032), .A2(n4608), .B1(n25033), .B2(n5328), .C1(
        n25034), .C2(n6240), .ZN(n25476) );
  OAI222D0 U8239 ( .A1(n25035), .A2(n6192), .B1(n25036), .B2(n4560), .C1(
        n25037), .C2(n5376), .ZN(n25475) );
  OAI22D0 U8240 ( .A1(n27079), .A2(n25038), .B1(n27078), .B2(n25039), .ZN(
        n25474) );
  OAI222D0 U8241 ( .A1(n24894), .A2(n25040), .B1(n25041), .B2(n5856), .C1(
        n25042), .C2(n5808), .ZN(n25473) );
  CKND0 U8242 ( .I(\Mem[44][10] ), .ZN(n24894) );
  AOI221D0 U8243 ( .A1(n27076), .A2(n25043), .B1(n27077), .B2(n25044), .C(
        n25477), .ZN(n25469) );
  OAI222D0 U8244 ( .A1(n25046), .A2(n6048), .B1(n24895), .B2(n25047), .C1(
        n25048), .C2(n4704), .ZN(n25477) );
  CKND0 U8245 ( .I(\Mem[45][10] ), .ZN(n24895) );
  NR4D0 U8246 ( .A1(n25478), .A2(n25479), .A3(n25480), .A4(n25481), .ZN(n25446) );
  OAI22D0 U8247 ( .A1(n25053), .A2(n5904), .B1(n25054), .B2(n5712), .ZN(n25481) );
  OAI222D0 U8248 ( .A1(n25055), .A2(n3840), .B1(n25056), .B2(n3888), .C1(
        n25057), .C2(n5952), .ZN(n25480) );
  OAI222D0 U8249 ( .A1(n25058), .A2(n3984), .B1(n25059), .B2(n4032), .C1(
        n25060), .C2(n3936), .ZN(n25479) );
  OAI222D0 U8250 ( .A1(n25061), .A2(n4128), .B1(n25062), .B2(n4176), .C1(
        n25063), .C2(n4080), .ZN(n25478) );
  NR4D0 U8251 ( .A1(n25482), .A2(n25483), .A3(n25484), .A4(n25485), .ZN(n25445) );
  OAI22D0 U8252 ( .A1(n25068), .A2(n2400), .B1(n25069), .B2(n2928), .ZN(n25485) );
  OAI222D0 U8253 ( .A1(n25070), .A2(n2496), .B1(n25071), .B2(n4320), .C1(
        n25072), .C2(n2640), .ZN(n25484) );
  OAI222D0 U8254 ( .A1(n25073), .A2(n4272), .B1(n24930), .B2(n3312), .C1(
        n25074), .C2(n4224), .ZN(n25483) );
  OAI222D0 U8255 ( .A1(n24932), .A2(n3408), .B1(n25075), .B2(n4848), .C1(
        n24931), .C2(n3360), .ZN(n25482) );
  ND4D0 U8256 ( .A1(n25486), .A2(n25487), .A3(n25488), .A4(n25489), .ZN(n2206)
         );
  AN4D0 U8257 ( .A1(n25490), .A2(n25491), .A3(n25492), .A4(n25493), .Z(n25489)
         );
  NR4D0 U8258 ( .A1(n25494), .A2(n25495), .A3(n25496), .A4(n25497), .ZN(n25493) );
  OAI222D0 U8259 ( .A1(n24979), .A2(n15493), .B1(n24980), .B2(n4463), .C1(
        n24964), .C2(n2255), .ZN(n25497) );
  OAI222D0 U8260 ( .A1(n24920), .A2(n2543), .B1(n24981), .B2(n5183), .C1(
        n24963), .C2(n2447), .ZN(n25496) );
  OAI222D0 U8261 ( .A1(n24982), .A2(n4943), .B1(n24983), .B2(n4991), .C1(
        n24984), .C2(n4895), .ZN(n25495) );
  OAI222D0 U8262 ( .A1(n24985), .A2(n4415), .B1(n24986), .B2(n3791), .C1(
        n24987), .C2(n4367), .ZN(n25494) );
  NR4D0 U8263 ( .A1(n25498), .A2(n25499), .A3(n25500), .A4(n25501), .ZN(n25492) );
  OAI22D0 U8264 ( .A1(n24922), .A2(n2831), .B1(n24992), .B2(n3743), .ZN(n25501) );
  OAI222D0 U8265 ( .A1(n24993), .A2(n17959), .B1(n24962), .B2(n2783), .C1(
        n24994), .C2(n17960), .ZN(n25500) );
  OAI222D0 U8266 ( .A1(n24995), .A2(n5231), .B1(n24961), .B2(n2687), .C1(
        n24921), .C2(n2735), .ZN(n25499) );
  OAI222D0 U8267 ( .A1(n24927), .A2(n3167), .B1(n24996), .B2(n4799), .C1(
        n24997), .C2(n15492), .ZN(n25498) );
  NR4D0 U8268 ( .A1(n25502), .A2(n25503), .A3(n25504), .A4(n25505), .ZN(n25491) );
  OAI22D0 U8269 ( .A1(n24928), .A2(n3215), .B1(n24926), .B2(n3119), .ZN(n25505) );
  OAI222D0 U8270 ( .A1(n25002), .A2(n3455), .B1(n24929), .B2(n3263), .C1(
        n24933), .C2(n2351), .ZN(n25504) );
  OAI222D0 U8271 ( .A1(n25003), .A2(n3599), .B1(n25004), .B2(n3503), .C1(
        n25005), .C2(n3551), .ZN(n25503) );
  OAI222D0 U8272 ( .A1(n24965), .A2(n2591), .B1(n25006), .B2(n3647), .C1(
        n25007), .C2(n3695), .ZN(n25502) );
  NR4D0 U8273 ( .A1(n25506), .A2(n25507), .A3(n25508), .A4(n25509), .ZN(n25490) );
  OAI22D0 U8274 ( .A1(n25012), .A2(n5135), .B1(n24966), .B2(n2303), .ZN(n25509) );
  OAI222D0 U8275 ( .A1(n24925), .A2(n3071), .B1(n24923), .B2(n2975), .C1(
        n24960), .C2(n2879), .ZN(n25508) );
  OAI222D0 U8276 ( .A1(n25013), .A2(n5519), .B1(n25014), .B2(n5567), .C1(
        n24924), .C2(n3023), .ZN(n25507) );
  OAI222D0 U8277 ( .A1(n25015), .A2(n6095), .B1(n25016), .B2(n5999), .C1(
        n25017), .C2(n6143), .ZN(n25506) );
  INR4D0 U8278 ( .A1(n25510), .B1(n25511), .B2(n25512), .B3(n25513), .ZN(
        n25488) );
  OAI222D0 U8279 ( .A1(n25022), .A2(n5471), .B1(n25023), .B2(n6335), .C1(
        n25024), .C2(n5423), .ZN(n25513) );
  OAI222D0 U8280 ( .A1(n25025), .A2(n4511), .B1(n25026), .B2(n24592), .C1(
        n25027), .C2(n5615), .ZN(n25512) );
  OR4D0 U8281 ( .A1(n25514), .A2(n25515), .A3(n25516), .A4(n25517), .Z(n25511)
         );
  OAI222D0 U8282 ( .A1(n25032), .A2(n4607), .B1(n25033), .B2(n5327), .C1(
        n25034), .C2(n6239), .ZN(n25517) );
  OAI222D0 U8283 ( .A1(n25035), .A2(n6191), .B1(n25036), .B2(n4559), .C1(
        n25037), .C2(n5375), .ZN(n25516) );
  OAI22D0 U8284 ( .A1(n27083), .A2(n25038), .B1(n27082), .B2(n25039), .ZN(
        n25515) );
  OAI222D0 U8285 ( .A1(n24892), .A2(n25040), .B1(n25041), .B2(n5855), .C1(
        n25042), .C2(n5807), .ZN(n25514) );
  CKND0 U8286 ( .I(\Mem[44][11] ), .ZN(n24892) );
  AOI221D0 U8287 ( .A1(n27080), .A2(n25043), .B1(n27081), .B2(n25044), .C(
        n25518), .ZN(n25510) );
  OAI222D0 U8288 ( .A1(n25046), .A2(n6047), .B1(n24893), .B2(n25047), .C1(
        n25048), .C2(n4703), .ZN(n25518) );
  CKND0 U8289 ( .I(\Mem[45][11] ), .ZN(n24893) );
  NR4D0 U8290 ( .A1(n25519), .A2(n25520), .A3(n25521), .A4(n25522), .ZN(n25487) );
  OAI22D0 U8291 ( .A1(n25053), .A2(n5903), .B1(n25054), .B2(n5711), .ZN(n25522) );
  OAI222D0 U8292 ( .A1(n25055), .A2(n3839), .B1(n25056), .B2(n3887), .C1(
        n25057), .C2(n5951), .ZN(n25521) );
  OAI222D0 U8293 ( .A1(n25058), .A2(n3983), .B1(n25059), .B2(n4031), .C1(
        n25060), .C2(n3935), .ZN(n25520) );
  OAI222D0 U8294 ( .A1(n25061), .A2(n4127), .B1(n25062), .B2(n4175), .C1(
        n25063), .C2(n4079), .ZN(n25519) );
  NR4D0 U8295 ( .A1(n25523), .A2(n25524), .A3(n25525), .A4(n25526), .ZN(n25486) );
  OAI22D0 U8296 ( .A1(n25068), .A2(n2399), .B1(n25069), .B2(n2927), .ZN(n25526) );
  OAI222D0 U8297 ( .A1(n25070), .A2(n2495), .B1(n25071), .B2(n4319), .C1(
        n25072), .C2(n2639), .ZN(n25525) );
  OAI222D0 U8298 ( .A1(n25073), .A2(n4271), .B1(n24930), .B2(n3311), .C1(
        n25074), .C2(n4223), .ZN(n25524) );
  OAI222D0 U8299 ( .A1(n24932), .A2(n3407), .B1(n25075), .B2(n4847), .C1(
        n24931), .C2(n3359), .ZN(n25523) );
  ND4D0 U8300 ( .A1(n25527), .A2(n25528), .A3(n25529), .A4(n25530), .ZN(n2205)
         );
  AN4D0 U8301 ( .A1(n25531), .A2(n25532), .A3(n25533), .A4(n25534), .Z(n25530)
         );
  NR4D0 U8302 ( .A1(n25535), .A2(n25536), .A3(n25537), .A4(n25538), .ZN(n25534) );
  OAI222D0 U8303 ( .A1(n24979), .A2(n15497), .B1(n24980), .B2(n4462), .C1(
        n24964), .C2(n2254), .ZN(n25538) );
  OAI222D0 U8304 ( .A1(n24920), .A2(n2542), .B1(n24981), .B2(n5182), .C1(
        n24963), .C2(n2446), .ZN(n25537) );
  OAI222D0 U8305 ( .A1(n24982), .A2(n4942), .B1(n24983), .B2(n4990), .C1(
        n24984), .C2(n4894), .ZN(n25536) );
  OAI222D0 U8306 ( .A1(n24985), .A2(n4414), .B1(n24986), .B2(n3790), .C1(
        n24987), .C2(n4366), .ZN(n25535) );
  NR4D0 U8307 ( .A1(n25539), .A2(n25540), .A3(n25541), .A4(n25542), .ZN(n25533) );
  OAI22D0 U8308 ( .A1(n24922), .A2(n2830), .B1(n24992), .B2(n3742), .ZN(n25542) );
  OAI222D0 U8309 ( .A1(n24993), .A2(n17962), .B1(n24962), .B2(n2782), .C1(
        n24994), .C2(n17963), .ZN(n25541) );
  OAI222D0 U8310 ( .A1(n24995), .A2(n5230), .B1(n24961), .B2(n2686), .C1(
        n24921), .C2(n2734), .ZN(n25540) );
  OAI222D0 U8311 ( .A1(n24927), .A2(n3166), .B1(n24996), .B2(n4798), .C1(
        n24997), .C2(n15496), .ZN(n25539) );
  NR4D0 U8312 ( .A1(n25543), .A2(n25544), .A3(n25545), .A4(n25546), .ZN(n25532) );
  OAI22D0 U8313 ( .A1(n24928), .A2(n3214), .B1(n24926), .B2(n3118), .ZN(n25546) );
  OAI222D0 U8314 ( .A1(n25002), .A2(n3454), .B1(n24929), .B2(n3262), .C1(
        n24933), .C2(n2350), .ZN(n25545) );
  OAI222D0 U8315 ( .A1(n25003), .A2(n3598), .B1(n25004), .B2(n3502), .C1(
        n25005), .C2(n3550), .ZN(n25544) );
  OAI222D0 U8316 ( .A1(n24965), .A2(n2590), .B1(n25006), .B2(n3646), .C1(
        n25007), .C2(n3694), .ZN(n25543) );
  NR4D0 U8317 ( .A1(n25547), .A2(n25548), .A3(n25549), .A4(n25550), .ZN(n25531) );
  OAI22D0 U8318 ( .A1(n25012), .A2(n5134), .B1(n24966), .B2(n2302), .ZN(n25550) );
  OAI222D0 U8319 ( .A1(n24925), .A2(n3070), .B1(n24923), .B2(n2974), .C1(
        n24960), .C2(n2878), .ZN(n25549) );
  OAI222D0 U8320 ( .A1(n25013), .A2(n5518), .B1(n25014), .B2(n5566), .C1(
        n24924), .C2(n3022), .ZN(n25548) );
  OAI222D0 U8321 ( .A1(n25015), .A2(n6094), .B1(n25016), .B2(n5998), .C1(
        n25017), .C2(n6142), .ZN(n25547) );
  INR4D0 U8322 ( .A1(n25551), .B1(n25552), .B2(n25553), .B3(n25554), .ZN(
        n25529) );
  OAI222D0 U8323 ( .A1(n25022), .A2(n5470), .B1(n25023), .B2(n6334), .C1(
        n25024), .C2(n5422), .ZN(n25554) );
  OAI222D0 U8324 ( .A1(n25025), .A2(n4510), .B1(n25026), .B2(n24595), .C1(
        n25027), .C2(n5614), .ZN(n25553) );
  OR4D0 U8325 ( .A1(n25555), .A2(n25556), .A3(n25557), .A4(n25558), .Z(n25552)
         );
  OAI222D0 U8326 ( .A1(n25032), .A2(n4606), .B1(n25033), .B2(n5326), .C1(
        n25034), .C2(n6238), .ZN(n25558) );
  OAI222D0 U8327 ( .A1(n25035), .A2(n6190), .B1(n25036), .B2(n4558), .C1(
        n25037), .C2(n5374), .ZN(n25557) );
  OAI22D0 U8328 ( .A1(n27087), .A2(n25038), .B1(n27086), .B2(n25039), .ZN(
        n25556) );
  OAI222D0 U8329 ( .A1(n24890), .A2(n25040), .B1(n25041), .B2(n5854), .C1(
        n25042), .C2(n5806), .ZN(n25555) );
  CKND0 U8330 ( .I(\Mem[44][12] ), .ZN(n24890) );
  AOI221D0 U8331 ( .A1(n27084), .A2(n25043), .B1(n27085), .B2(n25044), .C(
        n25559), .ZN(n25551) );
  OAI222D0 U8332 ( .A1(n25046), .A2(n6046), .B1(n24891), .B2(n25047), .C1(
        n25048), .C2(n4702), .ZN(n25559) );
  CKND0 U8333 ( .I(\Mem[45][12] ), .ZN(n24891) );
  NR4D0 U8334 ( .A1(n25560), .A2(n25561), .A3(n25562), .A4(n25563), .ZN(n25528) );
  OAI22D0 U8335 ( .A1(n25053), .A2(n5902), .B1(n25054), .B2(n5710), .ZN(n25563) );
  OAI222D0 U8336 ( .A1(n25055), .A2(n3838), .B1(n25056), .B2(n3886), .C1(
        n25057), .C2(n5950), .ZN(n25562) );
  OAI222D0 U8337 ( .A1(n25058), .A2(n3982), .B1(n25059), .B2(n4030), .C1(
        n25060), .C2(n3934), .ZN(n25561) );
  OAI222D0 U8338 ( .A1(n25061), .A2(n4126), .B1(n25062), .B2(n4174), .C1(
        n25063), .C2(n4078), .ZN(n25560) );
  NR4D0 U8339 ( .A1(n25564), .A2(n25565), .A3(n25566), .A4(n25567), .ZN(n25527) );
  OAI22D0 U8340 ( .A1(n25068), .A2(n2398), .B1(n25069), .B2(n2926), .ZN(n25567) );
  OAI222D0 U8341 ( .A1(n25070), .A2(n2494), .B1(n25071), .B2(n4318), .C1(
        n25072), .C2(n2638), .ZN(n25566) );
  OAI222D0 U8342 ( .A1(n25073), .A2(n4270), .B1(n24930), .B2(n3310), .C1(
        n25074), .C2(n4222), .ZN(n25565) );
  OAI222D0 U8343 ( .A1(n24932), .A2(n3406), .B1(n25075), .B2(n4846), .C1(
        n24931), .C2(n3358), .ZN(n25564) );
  ND4D0 U8344 ( .A1(n25568), .A2(n25569), .A3(n25570), .A4(n25571), .ZN(n2204)
         );
  AN4D0 U8345 ( .A1(n25572), .A2(n25573), .A3(n25574), .A4(n25575), .Z(n25571)
         );
  NR4D0 U8346 ( .A1(n25576), .A2(n25577), .A3(n25578), .A4(n25579), .ZN(n25575) );
  OAI222D0 U8347 ( .A1(n24979), .A2(n15501), .B1(n24980), .B2(n4461), .C1(
        n24964), .C2(n2253), .ZN(n25579) );
  OAI222D0 U8348 ( .A1(n24920), .A2(n2541), .B1(n24981), .B2(n5181), .C1(
        n24963), .C2(n2445), .ZN(n25578) );
  OAI222D0 U8349 ( .A1(n24982), .A2(n4941), .B1(n24983), .B2(n4989), .C1(
        n24984), .C2(n4893), .ZN(n25577) );
  OAI222D0 U8350 ( .A1(n24985), .A2(n4413), .B1(n24986), .B2(n3789), .C1(
        n24987), .C2(n4365), .ZN(n25576) );
  NR4D0 U8351 ( .A1(n25580), .A2(n25581), .A3(n25582), .A4(n25583), .ZN(n25574) );
  OAI22D0 U8352 ( .A1(n24922), .A2(n2829), .B1(n24992), .B2(n3741), .ZN(n25583) );
  OAI222D0 U8353 ( .A1(n24993), .A2(n17965), .B1(n24962), .B2(n2781), .C1(
        n24994), .C2(n17966), .ZN(n25582) );
  OAI222D0 U8354 ( .A1(n24995), .A2(n5229), .B1(n24961), .B2(n2685), .C1(
        n24921), .C2(n2733), .ZN(n25581) );
  OAI222D0 U8355 ( .A1(n24927), .A2(n3165), .B1(n24996), .B2(n4797), .C1(
        n24997), .C2(n15500), .ZN(n25580) );
  NR4D0 U8356 ( .A1(n25584), .A2(n25585), .A3(n25586), .A4(n25587), .ZN(n25573) );
  OAI22D0 U8357 ( .A1(n24928), .A2(n3213), .B1(n24926), .B2(n3117), .ZN(n25587) );
  OAI222D0 U8358 ( .A1(n25002), .A2(n3453), .B1(n24929), .B2(n3261), .C1(
        n24933), .C2(n2349), .ZN(n25586) );
  OAI222D0 U8359 ( .A1(n25003), .A2(n3597), .B1(n25004), .B2(n3501), .C1(
        n25005), .C2(n3549), .ZN(n25585) );
  OAI222D0 U8360 ( .A1(n24965), .A2(n2589), .B1(n25006), .B2(n3645), .C1(
        n25007), .C2(n3693), .ZN(n25584) );
  NR4D0 U8361 ( .A1(n25588), .A2(n25589), .A3(n25590), .A4(n25591), .ZN(n25572) );
  OAI22D0 U8362 ( .A1(n25012), .A2(n5133), .B1(n24966), .B2(n2301), .ZN(n25591) );
  OAI222D0 U8363 ( .A1(n24925), .A2(n3069), .B1(n24923), .B2(n2973), .C1(
        n24960), .C2(n2877), .ZN(n25590) );
  OAI222D0 U8364 ( .A1(n25013), .A2(n5517), .B1(n25014), .B2(n5565), .C1(
        n24924), .C2(n3021), .ZN(n25589) );
  OAI222D0 U8365 ( .A1(n25015), .A2(n6093), .B1(n25016), .B2(n5997), .C1(
        n25017), .C2(n6141), .ZN(n25588) );
  INR4D0 U8366 ( .A1(n25592), .B1(n25593), .B2(n25594), .B3(n25595), .ZN(
        n25570) );
  OAI222D0 U8367 ( .A1(n25022), .A2(n5469), .B1(n25023), .B2(n6333), .C1(
        n25024), .C2(n5421), .ZN(n25595) );
  OAI222D0 U8368 ( .A1(n25025), .A2(n4509), .B1(n25026), .B2(n24598), .C1(
        n25027), .C2(n5613), .ZN(n25594) );
  OR4D0 U8369 ( .A1(n25596), .A2(n25597), .A3(n25598), .A4(n25599), .Z(n25593)
         );
  OAI222D0 U8370 ( .A1(n25032), .A2(n4605), .B1(n25033), .B2(n5325), .C1(
        n25034), .C2(n6237), .ZN(n25599) );
  OAI222D0 U8371 ( .A1(n25035), .A2(n6189), .B1(n25036), .B2(n4557), .C1(
        n25037), .C2(n5373), .ZN(n25598) );
  OAI22D0 U8372 ( .A1(n27091), .A2(n25038), .B1(n27090), .B2(n25039), .ZN(
        n25597) );
  OAI222D0 U8373 ( .A1(n24888), .A2(n25040), .B1(n25041), .B2(n5853), .C1(
        n25042), .C2(n5805), .ZN(n25596) );
  CKND0 U8374 ( .I(\Mem[44][13] ), .ZN(n24888) );
  AOI221D0 U8375 ( .A1(n27088), .A2(n25043), .B1(n27089), .B2(n25044), .C(
        n25600), .ZN(n25592) );
  OAI222D0 U8376 ( .A1(n25046), .A2(n6045), .B1(n24889), .B2(n25047), .C1(
        n25048), .C2(n4701), .ZN(n25600) );
  CKND0 U8377 ( .I(\Mem[45][13] ), .ZN(n24889) );
  NR4D0 U8378 ( .A1(n25601), .A2(n25602), .A3(n25603), .A4(n25604), .ZN(n25569) );
  OAI22D0 U8379 ( .A1(n25053), .A2(n5901), .B1(n25054), .B2(n5709), .ZN(n25604) );
  OAI222D0 U8380 ( .A1(n25055), .A2(n3837), .B1(n25056), .B2(n3885), .C1(
        n25057), .C2(n5949), .ZN(n25603) );
  OAI222D0 U8381 ( .A1(n25058), .A2(n3981), .B1(n25059), .B2(n4029), .C1(
        n25060), .C2(n3933), .ZN(n25602) );
  OAI222D0 U8382 ( .A1(n25061), .A2(n4125), .B1(n25062), .B2(n4173), .C1(
        n25063), .C2(n4077), .ZN(n25601) );
  NR4D0 U8383 ( .A1(n25605), .A2(n25606), .A3(n25607), .A4(n25608), .ZN(n25568) );
  OAI22D0 U8384 ( .A1(n25068), .A2(n2397), .B1(n25069), .B2(n2925), .ZN(n25608) );
  OAI222D0 U8385 ( .A1(n25070), .A2(n2493), .B1(n25071), .B2(n4317), .C1(
        n25072), .C2(n2637), .ZN(n25607) );
  OAI222D0 U8386 ( .A1(n25073), .A2(n4269), .B1(n24930), .B2(n3309), .C1(
        n25074), .C2(n4221), .ZN(n25606) );
  OAI222D0 U8387 ( .A1(n24932), .A2(n3405), .B1(n25075), .B2(n4845), .C1(
        n24931), .C2(n3357), .ZN(n25605) );
  ND4D0 U8388 ( .A1(n25609), .A2(n25610), .A3(n25611), .A4(n25612), .ZN(n2203)
         );
  AN4D0 U8389 ( .A1(n25613), .A2(n25614), .A3(n25615), .A4(n25616), .Z(n25612)
         );
  NR4D0 U8390 ( .A1(n25617), .A2(n25618), .A3(n25619), .A4(n25620), .ZN(n25616) );
  OAI222D0 U8391 ( .A1(n24979), .A2(n15505), .B1(n24980), .B2(n4460), .C1(
        n24964), .C2(n2252), .ZN(n25620) );
  OAI222D0 U8392 ( .A1(n24920), .A2(n2540), .B1(n24981), .B2(n5180), .C1(
        n24963), .C2(n2444), .ZN(n25619) );
  OAI222D0 U8393 ( .A1(n24982), .A2(n4940), .B1(n24983), .B2(n4988), .C1(
        n24984), .C2(n4892), .ZN(n25618) );
  OAI222D0 U8394 ( .A1(n24985), .A2(n4412), .B1(n24986), .B2(n3788), .C1(
        n24987), .C2(n4364), .ZN(n25617) );
  NR4D0 U8395 ( .A1(n25621), .A2(n25622), .A3(n25623), .A4(n25624), .ZN(n25615) );
  OAI22D0 U8396 ( .A1(n24922), .A2(n2828), .B1(n24992), .B2(n3740), .ZN(n25624) );
  OAI222D0 U8397 ( .A1(n24993), .A2(n17968), .B1(n24962), .B2(n2780), .C1(
        n24994), .C2(n17969), .ZN(n25623) );
  OAI222D0 U8398 ( .A1(n24995), .A2(n5228), .B1(n24961), .B2(n2684), .C1(
        n24921), .C2(n2732), .ZN(n25622) );
  OAI222D0 U8399 ( .A1(n24927), .A2(n3164), .B1(n24996), .B2(n4796), .C1(
        n24997), .C2(n15504), .ZN(n25621) );
  NR4D0 U8400 ( .A1(n25625), .A2(n25626), .A3(n25627), .A4(n25628), .ZN(n25614) );
  OAI22D0 U8401 ( .A1(n24928), .A2(n3212), .B1(n24926), .B2(n3116), .ZN(n25628) );
  OAI222D0 U8402 ( .A1(n25002), .A2(n3452), .B1(n24929), .B2(n3260), .C1(
        n24933), .C2(n2348), .ZN(n25627) );
  OAI222D0 U8403 ( .A1(n25003), .A2(n3596), .B1(n25004), .B2(n3500), .C1(
        n25005), .C2(n3548), .ZN(n25626) );
  OAI222D0 U8404 ( .A1(n24965), .A2(n2588), .B1(n25006), .B2(n3644), .C1(
        n25007), .C2(n3692), .ZN(n25625) );
  NR4D0 U8405 ( .A1(n25629), .A2(n25630), .A3(n25631), .A4(n25632), .ZN(n25613) );
  OAI22D0 U8406 ( .A1(n25012), .A2(n5132), .B1(n24966), .B2(n2300), .ZN(n25632) );
  OAI222D0 U8407 ( .A1(n24925), .A2(n3068), .B1(n24923), .B2(n2972), .C1(
        n24960), .C2(n2876), .ZN(n25631) );
  OAI222D0 U8408 ( .A1(n25013), .A2(n5516), .B1(n25014), .B2(n5564), .C1(
        n24924), .C2(n3020), .ZN(n25630) );
  OAI222D0 U8409 ( .A1(n25015), .A2(n6092), .B1(n25016), .B2(n5996), .C1(
        n25017), .C2(n6140), .ZN(n25629) );
  INR4D0 U8410 ( .A1(n25633), .B1(n25634), .B2(n25635), .B3(n25636), .ZN(
        n25611) );
  OAI222D0 U8411 ( .A1(n25022), .A2(n5468), .B1(n25023), .B2(n6332), .C1(
        n25024), .C2(n5420), .ZN(n25636) );
  OAI222D0 U8412 ( .A1(n25025), .A2(n4508), .B1(n25026), .B2(n24601), .C1(
        n25027), .C2(n5612), .ZN(n25635) );
  OR4D0 U8413 ( .A1(n25637), .A2(n25638), .A3(n25639), .A4(n25640), .Z(n25634)
         );
  OAI222D0 U8414 ( .A1(n25032), .A2(n4604), .B1(n25033), .B2(n5324), .C1(
        n25034), .C2(n6236), .ZN(n25640) );
  OAI222D0 U8415 ( .A1(n25035), .A2(n6188), .B1(n25036), .B2(n4556), .C1(
        n25037), .C2(n5372), .ZN(n25639) );
  OAI22D0 U8416 ( .A1(n27095), .A2(n25038), .B1(n27094), .B2(n25039), .ZN(
        n25638) );
  OAI222D0 U8417 ( .A1(n24886), .A2(n25040), .B1(n25041), .B2(n5852), .C1(
        n25042), .C2(n5804), .ZN(n25637) );
  CKND0 U8418 ( .I(\Mem[44][14] ), .ZN(n24886) );
  AOI221D0 U8419 ( .A1(n27092), .A2(n25043), .B1(n27093), .B2(n25044), .C(
        n25641), .ZN(n25633) );
  OAI222D0 U8420 ( .A1(n25046), .A2(n6044), .B1(n24887), .B2(n25047), .C1(
        n25048), .C2(n4700), .ZN(n25641) );
  CKND0 U8421 ( .I(\Mem[45][14] ), .ZN(n24887) );
  NR4D0 U8422 ( .A1(n25642), .A2(n25643), .A3(n25644), .A4(n25645), .ZN(n25610) );
  OAI22D0 U8423 ( .A1(n25053), .A2(n5900), .B1(n25054), .B2(n5708), .ZN(n25645) );
  OAI222D0 U8424 ( .A1(n25055), .A2(n3836), .B1(n25056), .B2(n3884), .C1(
        n25057), .C2(n5948), .ZN(n25644) );
  OAI222D0 U8425 ( .A1(n25058), .A2(n3980), .B1(n25059), .B2(n4028), .C1(
        n25060), .C2(n3932), .ZN(n25643) );
  OAI222D0 U8426 ( .A1(n25061), .A2(n4124), .B1(n25062), .B2(n4172), .C1(
        n25063), .C2(n4076), .ZN(n25642) );
  NR4D0 U8427 ( .A1(n25646), .A2(n25647), .A3(n25648), .A4(n25649), .ZN(n25609) );
  OAI22D0 U8428 ( .A1(n25068), .A2(n2396), .B1(n25069), .B2(n2924), .ZN(n25649) );
  OAI222D0 U8429 ( .A1(n25070), .A2(n2492), .B1(n25071), .B2(n4316), .C1(
        n25072), .C2(n2636), .ZN(n25648) );
  OAI222D0 U8430 ( .A1(n25073), .A2(n4268), .B1(n24930), .B2(n3308), .C1(
        n25074), .C2(n4220), .ZN(n25647) );
  OAI222D0 U8431 ( .A1(n24932), .A2(n3404), .B1(n25075), .B2(n4844), .C1(
        n24931), .C2(n3356), .ZN(n25646) );
  ND4D0 U8432 ( .A1(n25650), .A2(n25651), .A3(n25652), .A4(n25653), .ZN(n2202)
         );
  AN4D0 U8433 ( .A1(n25654), .A2(n25655), .A3(n25656), .A4(n25657), .Z(n25653)
         );
  NR4D0 U8434 ( .A1(n25658), .A2(n25659), .A3(n25660), .A4(n25661), .ZN(n25657) );
  OAI222D0 U8435 ( .A1(n24979), .A2(n15509), .B1(n24980), .B2(n4459), .C1(
        n24964), .C2(n2251), .ZN(n25661) );
  OAI222D0 U8436 ( .A1(n24920), .A2(n2539), .B1(n24981), .B2(n5179), .C1(
        n24963), .C2(n2443), .ZN(n25660) );
  OAI222D0 U8437 ( .A1(n24982), .A2(n4939), .B1(n24983), .B2(n4987), .C1(
        n24984), .C2(n4891), .ZN(n25659) );
  OAI222D0 U8438 ( .A1(n24985), .A2(n4411), .B1(n24986), .B2(n3787), .C1(
        n24987), .C2(n4363), .ZN(n25658) );
  NR4D0 U8439 ( .A1(n25662), .A2(n25663), .A3(n25664), .A4(n25665), .ZN(n25656) );
  OAI22D0 U8440 ( .A1(n24922), .A2(n2827), .B1(n24992), .B2(n3739), .ZN(n25665) );
  OAI222D0 U8441 ( .A1(n24993), .A2(n17971), .B1(n24962), .B2(n2779), .C1(
        n24994), .C2(n17972), .ZN(n25664) );
  OAI222D0 U8442 ( .A1(n24995), .A2(n5227), .B1(n24961), .B2(n2683), .C1(
        n24921), .C2(n2731), .ZN(n25663) );
  OAI222D0 U8443 ( .A1(n24927), .A2(n3163), .B1(n24996), .B2(n4795), .C1(
        n24997), .C2(n15508), .ZN(n25662) );
  NR4D0 U8444 ( .A1(n25666), .A2(n25667), .A3(n25668), .A4(n25669), .ZN(n25655) );
  OAI22D0 U8445 ( .A1(n24928), .A2(n3211), .B1(n24926), .B2(n3115), .ZN(n25669) );
  OAI222D0 U8446 ( .A1(n25002), .A2(n3451), .B1(n24929), .B2(n3259), .C1(
        n24933), .C2(n2347), .ZN(n25668) );
  OAI222D0 U8447 ( .A1(n25003), .A2(n3595), .B1(n25004), .B2(n3499), .C1(
        n25005), .C2(n3547), .ZN(n25667) );
  OAI222D0 U8448 ( .A1(n24965), .A2(n2587), .B1(n25006), .B2(n3643), .C1(
        n25007), .C2(n3691), .ZN(n25666) );
  NR4D0 U8449 ( .A1(n25670), .A2(n25671), .A3(n25672), .A4(n25673), .ZN(n25654) );
  OAI22D0 U8450 ( .A1(n25012), .A2(n5131), .B1(n24966), .B2(n2299), .ZN(n25673) );
  OAI222D0 U8451 ( .A1(n24925), .A2(n3067), .B1(n24923), .B2(n2971), .C1(
        n24960), .C2(n2875), .ZN(n25672) );
  OAI222D0 U8452 ( .A1(n25013), .A2(n5515), .B1(n25014), .B2(n5563), .C1(
        n24924), .C2(n3019), .ZN(n25671) );
  OAI222D0 U8453 ( .A1(n25015), .A2(n6091), .B1(n25016), .B2(n5995), .C1(
        n25017), .C2(n6139), .ZN(n25670) );
  INR4D0 U8454 ( .A1(n25674), .B1(n25675), .B2(n25676), .B3(n25677), .ZN(
        n25652) );
  OAI222D0 U8455 ( .A1(n25022), .A2(n5467), .B1(n25023), .B2(n6331), .C1(
        n25024), .C2(n5419), .ZN(n25677) );
  OAI222D0 U8456 ( .A1(n25025), .A2(n4507), .B1(n25026), .B2(n24604), .C1(
        n25027), .C2(n5611), .ZN(n25676) );
  OR4D0 U8457 ( .A1(n25678), .A2(n25679), .A3(n25680), .A4(n25681), .Z(n25675)
         );
  OAI222D0 U8458 ( .A1(n25032), .A2(n4603), .B1(n25033), .B2(n5323), .C1(
        n25034), .C2(n6235), .ZN(n25681) );
  OAI222D0 U8459 ( .A1(n25035), .A2(n6187), .B1(n25036), .B2(n4555), .C1(
        n25037), .C2(n5371), .ZN(n25680) );
  OAI22D0 U8460 ( .A1(n27099), .A2(n25038), .B1(n27098), .B2(n25039), .ZN(
        n25679) );
  OAI222D0 U8461 ( .A1(n24884), .A2(n25040), .B1(n25041), .B2(n5851), .C1(
        n25042), .C2(n5803), .ZN(n25678) );
  CKND0 U8462 ( .I(\Mem[44][15] ), .ZN(n24884) );
  AOI221D0 U8463 ( .A1(n27096), .A2(n25043), .B1(n27097), .B2(n25044), .C(
        n25682), .ZN(n25674) );
  OAI222D0 U8464 ( .A1(n25046), .A2(n6043), .B1(n24885), .B2(n25047), .C1(
        n25048), .C2(n4699), .ZN(n25682) );
  CKND0 U8465 ( .I(\Mem[45][15] ), .ZN(n24885) );
  NR4D0 U8466 ( .A1(n25683), .A2(n25684), .A3(n25685), .A4(n25686), .ZN(n25651) );
  OAI22D0 U8467 ( .A1(n25053), .A2(n5899), .B1(n25054), .B2(n5707), .ZN(n25686) );
  OAI222D0 U8468 ( .A1(n25055), .A2(n3835), .B1(n25056), .B2(n3883), .C1(
        n25057), .C2(n5947), .ZN(n25685) );
  OAI222D0 U8469 ( .A1(n25058), .A2(n3979), .B1(n25059), .B2(n4027), .C1(
        n25060), .C2(n3931), .ZN(n25684) );
  OAI222D0 U8470 ( .A1(n25061), .A2(n4123), .B1(n25062), .B2(n4171), .C1(
        n25063), .C2(n4075), .ZN(n25683) );
  NR4D0 U8471 ( .A1(n25687), .A2(n25688), .A3(n25689), .A4(n25690), .ZN(n25650) );
  OAI22D0 U8472 ( .A1(n25068), .A2(n2395), .B1(n25069), .B2(n2923), .ZN(n25690) );
  OAI222D0 U8473 ( .A1(n25070), .A2(n2491), .B1(n25071), .B2(n4315), .C1(
        n25072), .C2(n2635), .ZN(n25689) );
  OAI222D0 U8474 ( .A1(n25073), .A2(n4267), .B1(n24930), .B2(n3307), .C1(
        n25074), .C2(n4219), .ZN(n25688) );
  OAI222D0 U8475 ( .A1(n24932), .A2(n3403), .B1(n25075), .B2(n4843), .C1(
        n24931), .C2(n3355), .ZN(n25687) );
  ND4D0 U8476 ( .A1(n25691), .A2(n25692), .A3(n25693), .A4(n25694), .ZN(n2201)
         );
  AN4D0 U8477 ( .A1(n25695), .A2(n25696), .A3(n25697), .A4(n25698), .Z(n25694)
         );
  NR4D0 U8478 ( .A1(n25699), .A2(n25700), .A3(n25701), .A4(n25702), .ZN(n25698) );
  OAI222D0 U8479 ( .A1(n24979), .A2(n15513), .B1(n24980), .B2(n4458), .C1(
        n24964), .C2(n2250), .ZN(n25702) );
  OAI222D0 U8480 ( .A1(n24920), .A2(n2538), .B1(n24981), .B2(n5178), .C1(
        n24963), .C2(n2442), .ZN(n25701) );
  OAI222D0 U8481 ( .A1(n24982), .A2(n4938), .B1(n24983), .B2(n4986), .C1(
        n24984), .C2(n4890), .ZN(n25700) );
  OAI222D0 U8482 ( .A1(n24985), .A2(n4410), .B1(n24986), .B2(n3786), .C1(
        n24987), .C2(n4362), .ZN(n25699) );
  NR4D0 U8483 ( .A1(n25703), .A2(n25704), .A3(n25705), .A4(n25706), .ZN(n25697) );
  OAI22D0 U8484 ( .A1(n24922), .A2(n2826), .B1(n24992), .B2(n3738), .ZN(n25706) );
  OAI222D0 U8485 ( .A1(n24993), .A2(n17974), .B1(n24962), .B2(n2778), .C1(
        n24994), .C2(n17975), .ZN(n25705) );
  OAI222D0 U8486 ( .A1(n24995), .A2(n5226), .B1(n24961), .B2(n2682), .C1(
        n24921), .C2(n2730), .ZN(n25704) );
  OAI222D0 U8487 ( .A1(n24927), .A2(n3162), .B1(n24996), .B2(n4794), .C1(
        n24997), .C2(n15512), .ZN(n25703) );
  NR4D0 U8488 ( .A1(n25707), .A2(n25708), .A3(n25709), .A4(n25710), .ZN(n25696) );
  OAI22D0 U8489 ( .A1(n24928), .A2(n3210), .B1(n24926), .B2(n3114), .ZN(n25710) );
  OAI222D0 U8490 ( .A1(n25002), .A2(n3450), .B1(n24929), .B2(n3258), .C1(
        n24933), .C2(n2346), .ZN(n25709) );
  OAI222D0 U8491 ( .A1(n25003), .A2(n3594), .B1(n25004), .B2(n3498), .C1(
        n25005), .C2(n3546), .ZN(n25708) );
  OAI222D0 U8492 ( .A1(n24965), .A2(n2586), .B1(n25006), .B2(n3642), .C1(
        n25007), .C2(n3690), .ZN(n25707) );
  NR4D0 U8493 ( .A1(n25711), .A2(n25712), .A3(n25713), .A4(n25714), .ZN(n25695) );
  OAI22D0 U8494 ( .A1(n25012), .A2(n5130), .B1(n24966), .B2(n2298), .ZN(n25714) );
  OAI222D0 U8495 ( .A1(n24925), .A2(n3066), .B1(n24923), .B2(n2970), .C1(
        n24960), .C2(n2874), .ZN(n25713) );
  OAI222D0 U8496 ( .A1(n25013), .A2(n5514), .B1(n25014), .B2(n5562), .C1(
        n24924), .C2(n3018), .ZN(n25712) );
  OAI222D0 U8497 ( .A1(n25015), .A2(n6090), .B1(n25016), .B2(n5994), .C1(
        n25017), .C2(n6138), .ZN(n25711) );
  INR4D0 U8498 ( .A1(n25715), .B1(n25716), .B2(n25717), .B3(n25718), .ZN(
        n25693) );
  OAI222D0 U8499 ( .A1(n25022), .A2(n5466), .B1(n25023), .B2(n6330), .C1(
        n25024), .C2(n5418), .ZN(n25718) );
  OAI222D0 U8500 ( .A1(n25025), .A2(n4506), .B1(n25026), .B2(n24607), .C1(
        n25027), .C2(n5610), .ZN(n25717) );
  OR4D0 U8501 ( .A1(n25719), .A2(n25720), .A3(n25721), .A4(n25722), .Z(n25716)
         );
  OAI222D0 U8502 ( .A1(n25032), .A2(n4602), .B1(n25033), .B2(n5322), .C1(
        n25034), .C2(n6234), .ZN(n25722) );
  OAI222D0 U8503 ( .A1(n25035), .A2(n6186), .B1(n25036), .B2(n4554), .C1(
        n25037), .C2(n5370), .ZN(n25721) );
  OAI22D0 U8504 ( .A1(n27103), .A2(n25038), .B1(n27102), .B2(n25039), .ZN(
        n25720) );
  OAI222D0 U8505 ( .A1(n24882), .A2(n25040), .B1(n25041), .B2(n5850), .C1(
        n25042), .C2(n5802), .ZN(n25719) );
  CKND0 U8506 ( .I(\Mem[44][16] ), .ZN(n24882) );
  AOI221D0 U8507 ( .A1(n27100), .A2(n25043), .B1(n27101), .B2(n25044), .C(
        n25723), .ZN(n25715) );
  OAI222D0 U8508 ( .A1(n25046), .A2(n6042), .B1(n24883), .B2(n25047), .C1(
        n25048), .C2(n4698), .ZN(n25723) );
  CKND0 U8509 ( .I(\Mem[45][16] ), .ZN(n24883) );
  NR4D0 U8510 ( .A1(n25724), .A2(n25725), .A3(n25726), .A4(n25727), .ZN(n25692) );
  OAI22D0 U8511 ( .A1(n25053), .A2(n5898), .B1(n25054), .B2(n5706), .ZN(n25727) );
  OAI222D0 U8512 ( .A1(n25055), .A2(n3834), .B1(n25056), .B2(n3882), .C1(
        n25057), .C2(n5946), .ZN(n25726) );
  OAI222D0 U8513 ( .A1(n25058), .A2(n3978), .B1(n25059), .B2(n4026), .C1(
        n25060), .C2(n3930), .ZN(n25725) );
  OAI222D0 U8514 ( .A1(n25061), .A2(n4122), .B1(n25062), .B2(n4170), .C1(
        n25063), .C2(n4074), .ZN(n25724) );
  NR4D0 U8515 ( .A1(n25728), .A2(n25729), .A3(n25730), .A4(n25731), .ZN(n25691) );
  OAI22D0 U8516 ( .A1(n25068), .A2(n2394), .B1(n25069), .B2(n2922), .ZN(n25731) );
  OAI222D0 U8517 ( .A1(n25070), .A2(n2490), .B1(n25071), .B2(n4314), .C1(
        n25072), .C2(n2634), .ZN(n25730) );
  OAI222D0 U8518 ( .A1(n25073), .A2(n4266), .B1(n24930), .B2(n3306), .C1(
        n25074), .C2(n4218), .ZN(n25729) );
  OAI222D0 U8519 ( .A1(n24932), .A2(n3402), .B1(n25075), .B2(n4842), .C1(
        n24931), .C2(n3354), .ZN(n25728) );
  ND4D0 U8520 ( .A1(n25732), .A2(n25733), .A3(n25734), .A4(n25735), .ZN(n2200)
         );
  AN4D0 U8521 ( .A1(n25736), .A2(n25737), .A3(n25738), .A4(n25739), .Z(n25735)
         );
  NR4D0 U8522 ( .A1(n25740), .A2(n25741), .A3(n25742), .A4(n25743), .ZN(n25739) );
  OAI222D0 U8523 ( .A1(n24979), .A2(n15517), .B1(n24980), .B2(n4457), .C1(
        n24964), .C2(n2249), .ZN(n25743) );
  OAI222D0 U8524 ( .A1(n24920), .A2(n2537), .B1(n24981), .B2(n5177), .C1(
        n24963), .C2(n2441), .ZN(n25742) );
  OAI222D0 U8525 ( .A1(n24982), .A2(n4937), .B1(n24983), .B2(n4985), .C1(
        n24984), .C2(n4889), .ZN(n25741) );
  OAI222D0 U8526 ( .A1(n24985), .A2(n4409), .B1(n24986), .B2(n3785), .C1(
        n24987), .C2(n4361), .ZN(n25740) );
  NR4D0 U8527 ( .A1(n25744), .A2(n25745), .A3(n25746), .A4(n25747), .ZN(n25738) );
  OAI22D0 U8528 ( .A1(n24922), .A2(n2825), .B1(n24992), .B2(n3737), .ZN(n25747) );
  OAI222D0 U8529 ( .A1(n24993), .A2(n17977), .B1(n24962), .B2(n2777), .C1(
        n24994), .C2(n17978), .ZN(n25746) );
  OAI222D0 U8530 ( .A1(n24995), .A2(n5225), .B1(n24961), .B2(n2681), .C1(
        n24921), .C2(n2729), .ZN(n25745) );
  OAI222D0 U8531 ( .A1(n24927), .A2(n3161), .B1(n24996), .B2(n4793), .C1(
        n24997), .C2(n15516), .ZN(n25744) );
  NR4D0 U8532 ( .A1(n25748), .A2(n25749), .A3(n25750), .A4(n25751), .ZN(n25737) );
  OAI22D0 U8533 ( .A1(n24928), .A2(n3209), .B1(n24926), .B2(n3113), .ZN(n25751) );
  OAI222D0 U8534 ( .A1(n25002), .A2(n3449), .B1(n24929), .B2(n3257), .C1(
        n24933), .C2(n2345), .ZN(n25750) );
  OAI222D0 U8535 ( .A1(n25003), .A2(n3593), .B1(n25004), .B2(n3497), .C1(
        n25005), .C2(n3545), .ZN(n25749) );
  OAI222D0 U8536 ( .A1(n24965), .A2(n2585), .B1(n25006), .B2(n3641), .C1(
        n25007), .C2(n3689), .ZN(n25748) );
  NR4D0 U8537 ( .A1(n25752), .A2(n25753), .A3(n25754), .A4(n25755), .ZN(n25736) );
  OAI22D0 U8538 ( .A1(n25012), .A2(n5129), .B1(n24966), .B2(n2297), .ZN(n25755) );
  OAI222D0 U8539 ( .A1(n24925), .A2(n3065), .B1(n24923), .B2(n2969), .C1(
        n24960), .C2(n2873), .ZN(n25754) );
  OAI222D0 U8540 ( .A1(n25013), .A2(n5513), .B1(n25014), .B2(n5561), .C1(
        n24924), .C2(n3017), .ZN(n25753) );
  OAI222D0 U8541 ( .A1(n25015), .A2(n6089), .B1(n25016), .B2(n5993), .C1(
        n25017), .C2(n6137), .ZN(n25752) );
  INR4D0 U8542 ( .A1(n25756), .B1(n25757), .B2(n25758), .B3(n25759), .ZN(
        n25734) );
  OAI222D0 U8543 ( .A1(n25022), .A2(n5465), .B1(n25023), .B2(n6329), .C1(
        n25024), .C2(n5417), .ZN(n25759) );
  OAI222D0 U8544 ( .A1(n25025), .A2(n4505), .B1(n25026), .B2(n24610), .C1(
        n25027), .C2(n5609), .ZN(n25758) );
  OR4D0 U8545 ( .A1(n25760), .A2(n25761), .A3(n25762), .A4(n25763), .Z(n25757)
         );
  OAI222D0 U8546 ( .A1(n25032), .A2(n4601), .B1(n25033), .B2(n5321), .C1(
        n25034), .C2(n6233), .ZN(n25763) );
  OAI222D0 U8547 ( .A1(n25035), .A2(n6185), .B1(n25036), .B2(n4553), .C1(
        n25037), .C2(n5369), .ZN(n25762) );
  OAI22D0 U8548 ( .A1(n27107), .A2(n25038), .B1(n27106), .B2(n25039), .ZN(
        n25761) );
  OAI222D0 U8549 ( .A1(n24880), .A2(n25040), .B1(n25041), .B2(n5849), .C1(
        n25042), .C2(n5801), .ZN(n25760) );
  CKND0 U8550 ( .I(\Mem[44][17] ), .ZN(n24880) );
  AOI221D0 U8551 ( .A1(n27104), .A2(n25043), .B1(n27105), .B2(n25044), .C(
        n25764), .ZN(n25756) );
  OAI222D0 U8552 ( .A1(n25046), .A2(n6041), .B1(n24881), .B2(n25047), .C1(
        n25048), .C2(n4697), .ZN(n25764) );
  CKND0 U8553 ( .I(\Mem[45][17] ), .ZN(n24881) );
  NR4D0 U8554 ( .A1(n25765), .A2(n25766), .A3(n25767), .A4(n25768), .ZN(n25733) );
  OAI22D0 U8555 ( .A1(n25053), .A2(n5897), .B1(n25054), .B2(n5705), .ZN(n25768) );
  OAI222D0 U8556 ( .A1(n25055), .A2(n3833), .B1(n25056), .B2(n3881), .C1(
        n25057), .C2(n5945), .ZN(n25767) );
  OAI222D0 U8557 ( .A1(n25058), .A2(n3977), .B1(n25059), .B2(n4025), .C1(
        n25060), .C2(n3929), .ZN(n25766) );
  OAI222D0 U8558 ( .A1(n25061), .A2(n4121), .B1(n25062), .B2(n4169), .C1(
        n25063), .C2(n4073), .ZN(n25765) );
  NR4D0 U8559 ( .A1(n25769), .A2(n25770), .A3(n25771), .A4(n25772), .ZN(n25732) );
  OAI22D0 U8560 ( .A1(n25068), .A2(n2393), .B1(n25069), .B2(n2921), .ZN(n25772) );
  OAI222D0 U8561 ( .A1(n25070), .A2(n2489), .B1(n25071), .B2(n4313), .C1(
        n25072), .C2(n2633), .ZN(n25771) );
  OAI222D0 U8562 ( .A1(n25073), .A2(n4265), .B1(n24930), .B2(n3305), .C1(
        n25074), .C2(n4217), .ZN(n25770) );
  OAI222D0 U8563 ( .A1(n24932), .A2(n3401), .B1(n25075), .B2(n4841), .C1(
        n24931), .C2(n3353), .ZN(n25769) );
  ND4D0 U8564 ( .A1(n25773), .A2(n25774), .A3(n25775), .A4(n25776), .ZN(n2199)
         );
  AN4D0 U8565 ( .A1(n25777), .A2(n25778), .A3(n25779), .A4(n25780), .Z(n25776)
         );
  NR4D0 U8566 ( .A1(n25781), .A2(n25782), .A3(n25783), .A4(n25784), .ZN(n25780) );
  OAI222D0 U8567 ( .A1(n24979), .A2(n15521), .B1(n24980), .B2(n4456), .C1(
        n24964), .C2(n2248), .ZN(n25784) );
  OAI222D0 U8568 ( .A1(n24920), .A2(n2536), .B1(n24981), .B2(n5176), .C1(
        n24963), .C2(n2440), .ZN(n25783) );
  OAI222D0 U8569 ( .A1(n24982), .A2(n4936), .B1(n24983), .B2(n4984), .C1(
        n24984), .C2(n4888), .ZN(n25782) );
  OAI222D0 U8570 ( .A1(n24985), .A2(n4408), .B1(n24986), .B2(n3784), .C1(
        n24987), .C2(n4360), .ZN(n25781) );
  NR4D0 U8571 ( .A1(n25785), .A2(n25786), .A3(n25787), .A4(n25788), .ZN(n25779) );
  OAI22D0 U8572 ( .A1(n24922), .A2(n2824), .B1(n24992), .B2(n3736), .ZN(n25788) );
  OAI222D0 U8573 ( .A1(n24993), .A2(n17980), .B1(n24962), .B2(n2776), .C1(
        n24994), .C2(n17981), .ZN(n25787) );
  OAI222D0 U8574 ( .A1(n24995), .A2(n5224), .B1(n24961), .B2(n2680), .C1(
        n24921), .C2(n2728), .ZN(n25786) );
  OAI222D0 U8575 ( .A1(n24927), .A2(n3160), .B1(n24996), .B2(n4792), .C1(
        n24997), .C2(n15520), .ZN(n25785) );
  NR4D0 U8576 ( .A1(n25789), .A2(n25790), .A3(n25791), .A4(n25792), .ZN(n25778) );
  OAI22D0 U8577 ( .A1(n24928), .A2(n3208), .B1(n24926), .B2(n3112), .ZN(n25792) );
  OAI222D0 U8578 ( .A1(n25002), .A2(n3448), .B1(n24929), .B2(n3256), .C1(
        n24933), .C2(n2344), .ZN(n25791) );
  OAI222D0 U8579 ( .A1(n25003), .A2(n3592), .B1(n25004), .B2(n3496), .C1(
        n25005), .C2(n3544), .ZN(n25790) );
  OAI222D0 U8580 ( .A1(n24965), .A2(n2584), .B1(n25006), .B2(n3640), .C1(
        n25007), .C2(n3688), .ZN(n25789) );
  NR4D0 U8581 ( .A1(n25793), .A2(n25794), .A3(n25795), .A4(n25796), .ZN(n25777) );
  OAI22D0 U8582 ( .A1(n25012), .A2(n5128), .B1(n24966), .B2(n2296), .ZN(n25796) );
  OAI222D0 U8583 ( .A1(n24925), .A2(n3064), .B1(n24923), .B2(n2968), .C1(
        n24960), .C2(n2872), .ZN(n25795) );
  OAI222D0 U8584 ( .A1(n25013), .A2(n5512), .B1(n25014), .B2(n5560), .C1(
        n24924), .C2(n3016), .ZN(n25794) );
  OAI222D0 U8585 ( .A1(n25015), .A2(n6088), .B1(n25016), .B2(n5992), .C1(
        n25017), .C2(n6136), .ZN(n25793) );
  INR4D0 U8586 ( .A1(n25797), .B1(n25798), .B2(n25799), .B3(n25800), .ZN(
        n25775) );
  OAI222D0 U8587 ( .A1(n25022), .A2(n5464), .B1(n25023), .B2(n6328), .C1(
        n25024), .C2(n5416), .ZN(n25800) );
  OAI222D0 U8588 ( .A1(n25025), .A2(n4504), .B1(n25026), .B2(n24613), .C1(
        n25027), .C2(n5608), .ZN(n25799) );
  OR4D0 U8589 ( .A1(n25801), .A2(n25802), .A3(n25803), .A4(n25804), .Z(n25798)
         );
  OAI222D0 U8590 ( .A1(n25032), .A2(n4600), .B1(n25033), .B2(n5320), .C1(
        n25034), .C2(n6232), .ZN(n25804) );
  OAI222D0 U8591 ( .A1(n25035), .A2(n6184), .B1(n25036), .B2(n4552), .C1(
        n25037), .C2(n5368), .ZN(n25803) );
  OAI22D0 U8592 ( .A1(n27111), .A2(n25038), .B1(n27110), .B2(n25039), .ZN(
        n25802) );
  OAI222D0 U8593 ( .A1(n24878), .A2(n25040), .B1(n25041), .B2(n5848), .C1(
        n25042), .C2(n5800), .ZN(n25801) );
  CKND0 U8594 ( .I(\Mem[44][18] ), .ZN(n24878) );
  AOI221D0 U8595 ( .A1(n27108), .A2(n25043), .B1(n27109), .B2(n25044), .C(
        n25805), .ZN(n25797) );
  OAI222D0 U8596 ( .A1(n25046), .A2(n6040), .B1(n24879), .B2(n25047), .C1(
        n25048), .C2(n4696), .ZN(n25805) );
  CKND0 U8597 ( .I(\Mem[45][18] ), .ZN(n24879) );
  NR4D0 U8598 ( .A1(n25806), .A2(n25807), .A3(n25808), .A4(n25809), .ZN(n25774) );
  OAI22D0 U8599 ( .A1(n25053), .A2(n5896), .B1(n25054), .B2(n5704), .ZN(n25809) );
  OAI222D0 U8600 ( .A1(n25055), .A2(n3832), .B1(n25056), .B2(n3880), .C1(
        n25057), .C2(n5944), .ZN(n25808) );
  OAI222D0 U8601 ( .A1(n25058), .A2(n3976), .B1(n25059), .B2(n4024), .C1(
        n25060), .C2(n3928), .ZN(n25807) );
  OAI222D0 U8602 ( .A1(n25061), .A2(n4120), .B1(n25062), .B2(n4168), .C1(
        n25063), .C2(n4072), .ZN(n25806) );
  NR4D0 U8603 ( .A1(n25810), .A2(n25811), .A3(n25812), .A4(n25813), .ZN(n25773) );
  OAI22D0 U8604 ( .A1(n25068), .A2(n2392), .B1(n25069), .B2(n2920), .ZN(n25813) );
  OAI222D0 U8605 ( .A1(n25070), .A2(n2488), .B1(n25071), .B2(n4312), .C1(
        n25072), .C2(n2632), .ZN(n25812) );
  OAI222D0 U8606 ( .A1(n25073), .A2(n4264), .B1(n24930), .B2(n3304), .C1(
        n25074), .C2(n4216), .ZN(n25811) );
  OAI222D0 U8607 ( .A1(n24932), .A2(n3400), .B1(n25075), .B2(n4840), .C1(
        n24931), .C2(n3352), .ZN(n25810) );
  ND4D0 U8608 ( .A1(n25814), .A2(n25815), .A3(n25816), .A4(n25817), .ZN(n2198)
         );
  AN4D0 U8609 ( .A1(n25818), .A2(n25819), .A3(n25820), .A4(n25821), .Z(n25817)
         );
  NR4D0 U8610 ( .A1(n25822), .A2(n25823), .A3(n25824), .A4(n25825), .ZN(n25821) );
  OAI222D0 U8611 ( .A1(n24979), .A2(n15525), .B1(n24980), .B2(n4455), .C1(
        n24964), .C2(n2247), .ZN(n25825) );
  OAI222D0 U8612 ( .A1(n24920), .A2(n2535), .B1(n24981), .B2(n5175), .C1(
        n24963), .C2(n2439), .ZN(n25824) );
  OAI222D0 U8613 ( .A1(n24982), .A2(n4935), .B1(n24983), .B2(n4983), .C1(
        n24984), .C2(n4887), .ZN(n25823) );
  OAI222D0 U8614 ( .A1(n24985), .A2(n4407), .B1(n24986), .B2(n3783), .C1(
        n24987), .C2(n4359), .ZN(n25822) );
  NR4D0 U8615 ( .A1(n25826), .A2(n25827), .A3(n25828), .A4(n25829), .ZN(n25820) );
  OAI22D0 U8616 ( .A1(n24922), .A2(n2823), .B1(n24992), .B2(n3735), .ZN(n25829) );
  OAI222D0 U8617 ( .A1(n24993), .A2(n17983), .B1(n24962), .B2(n2775), .C1(
        n24994), .C2(n17984), .ZN(n25828) );
  OAI222D0 U8618 ( .A1(n24995), .A2(n5223), .B1(n24961), .B2(n2679), .C1(
        n24921), .C2(n2727), .ZN(n25827) );
  OAI222D0 U8619 ( .A1(n24927), .A2(n3159), .B1(n24996), .B2(n4791), .C1(
        n24997), .C2(n15524), .ZN(n25826) );
  NR4D0 U8620 ( .A1(n25830), .A2(n25831), .A3(n25832), .A4(n25833), .ZN(n25819) );
  OAI22D0 U8621 ( .A1(n24928), .A2(n3207), .B1(n24926), .B2(n3111), .ZN(n25833) );
  OAI222D0 U8622 ( .A1(n25002), .A2(n3447), .B1(n24929), .B2(n3255), .C1(
        n24933), .C2(n2343), .ZN(n25832) );
  OAI222D0 U8623 ( .A1(n25003), .A2(n3591), .B1(n25004), .B2(n3495), .C1(
        n25005), .C2(n3543), .ZN(n25831) );
  OAI222D0 U8624 ( .A1(n24965), .A2(n2583), .B1(n25006), .B2(n3639), .C1(
        n25007), .C2(n3687), .ZN(n25830) );
  NR4D0 U8625 ( .A1(n25834), .A2(n25835), .A3(n25836), .A4(n25837), .ZN(n25818) );
  OAI22D0 U8626 ( .A1(n25012), .A2(n5127), .B1(n24966), .B2(n2295), .ZN(n25837) );
  OAI222D0 U8627 ( .A1(n24925), .A2(n3063), .B1(n24923), .B2(n2967), .C1(
        n24960), .C2(n2871), .ZN(n25836) );
  OAI222D0 U8628 ( .A1(n25013), .A2(n5511), .B1(n25014), .B2(n5559), .C1(
        n24924), .C2(n3015), .ZN(n25835) );
  OAI222D0 U8629 ( .A1(n25015), .A2(n6087), .B1(n25016), .B2(n5991), .C1(
        n25017), .C2(n6135), .ZN(n25834) );
  INR4D0 U8630 ( .A1(n25838), .B1(n25839), .B2(n25840), .B3(n25841), .ZN(
        n25816) );
  OAI222D0 U8631 ( .A1(n25022), .A2(n5463), .B1(n25023), .B2(n6327), .C1(
        n25024), .C2(n5415), .ZN(n25841) );
  OAI222D0 U8632 ( .A1(n25025), .A2(n4503), .B1(n25026), .B2(n24616), .C1(
        n25027), .C2(n5607), .ZN(n25840) );
  OR4D0 U8633 ( .A1(n25842), .A2(n25843), .A3(n25844), .A4(n25845), .Z(n25839)
         );
  OAI222D0 U8634 ( .A1(n25032), .A2(n4599), .B1(n25033), .B2(n5319), .C1(
        n25034), .C2(n6231), .ZN(n25845) );
  OAI222D0 U8635 ( .A1(n25035), .A2(n6183), .B1(n25036), .B2(n4551), .C1(
        n25037), .C2(n5367), .ZN(n25844) );
  OAI22D0 U8636 ( .A1(n27115), .A2(n25038), .B1(n27114), .B2(n25039), .ZN(
        n25843) );
  OAI222D0 U8637 ( .A1(n24876), .A2(n25040), .B1(n25041), .B2(n5847), .C1(
        n25042), .C2(n5799), .ZN(n25842) );
  CKND0 U8638 ( .I(\Mem[44][19] ), .ZN(n24876) );
  AOI221D0 U8639 ( .A1(n27112), .A2(n25043), .B1(n27113), .B2(n25044), .C(
        n25846), .ZN(n25838) );
  OAI222D0 U8640 ( .A1(n25046), .A2(n6039), .B1(n24877), .B2(n25047), .C1(
        n25048), .C2(n4695), .ZN(n25846) );
  CKND0 U8641 ( .I(\Mem[45][19] ), .ZN(n24877) );
  NR4D0 U8642 ( .A1(n25847), .A2(n25848), .A3(n25849), .A4(n25850), .ZN(n25815) );
  OAI22D0 U8643 ( .A1(n25053), .A2(n5895), .B1(n25054), .B2(n5703), .ZN(n25850) );
  OAI222D0 U8644 ( .A1(n25055), .A2(n3831), .B1(n25056), .B2(n3879), .C1(
        n25057), .C2(n5943), .ZN(n25849) );
  OAI222D0 U8645 ( .A1(n25058), .A2(n3975), .B1(n25059), .B2(n4023), .C1(
        n25060), .C2(n3927), .ZN(n25848) );
  OAI222D0 U8646 ( .A1(n25061), .A2(n4119), .B1(n25062), .B2(n4167), .C1(
        n25063), .C2(n4071), .ZN(n25847) );
  NR4D0 U8647 ( .A1(n25851), .A2(n25852), .A3(n25853), .A4(n25854), .ZN(n25814) );
  OAI22D0 U8648 ( .A1(n25068), .A2(n2391), .B1(n25069), .B2(n2919), .ZN(n25854) );
  OAI222D0 U8649 ( .A1(n25070), .A2(n2487), .B1(n25071), .B2(n4311), .C1(
        n25072), .C2(n2631), .ZN(n25853) );
  OAI222D0 U8650 ( .A1(n25073), .A2(n4263), .B1(n24930), .B2(n3303), .C1(
        n25074), .C2(n4215), .ZN(n25852) );
  OAI222D0 U8651 ( .A1(n24932), .A2(n3399), .B1(n25075), .B2(n4839), .C1(
        n24931), .C2(n3351), .ZN(n25851) );
  ND4D0 U8652 ( .A1(n25855), .A2(n25856), .A3(n25857), .A4(n25858), .ZN(n2197)
         );
  AN4D0 U8653 ( .A1(n25859), .A2(n25860), .A3(n25861), .A4(n25862), .Z(n25858)
         );
  NR4D0 U8654 ( .A1(n25863), .A2(n25864), .A3(n25865), .A4(n25866), .ZN(n25862) );
  OAI222D0 U8655 ( .A1(n24979), .A2(n15529), .B1(n24980), .B2(n4454), .C1(
        n24964), .C2(n2246), .ZN(n25866) );
  OAI222D0 U8656 ( .A1(n24920), .A2(n2534), .B1(n24981), .B2(n5174), .C1(
        n24963), .C2(n2438), .ZN(n25865) );
  OAI222D0 U8657 ( .A1(n24982), .A2(n4934), .B1(n24983), .B2(n4982), .C1(
        n24984), .C2(n4886), .ZN(n25864) );
  OAI222D0 U8658 ( .A1(n24985), .A2(n4406), .B1(n24986), .B2(n3782), .C1(
        n24987), .C2(n4358), .ZN(n25863) );
  NR4D0 U8659 ( .A1(n25867), .A2(n25868), .A3(n25869), .A4(n25870), .ZN(n25861) );
  OAI22D0 U8660 ( .A1(n24922), .A2(n2822), .B1(n24992), .B2(n3734), .ZN(n25870) );
  OAI222D0 U8661 ( .A1(n24993), .A2(n17986), .B1(n24962), .B2(n2774), .C1(
        n24994), .C2(n17987), .ZN(n25869) );
  OAI222D0 U8662 ( .A1(n24995), .A2(n5222), .B1(n24961), .B2(n2678), .C1(
        n24921), .C2(n2726), .ZN(n25868) );
  OAI222D0 U8663 ( .A1(n24927), .A2(n3158), .B1(n24996), .B2(n4790), .C1(
        n24997), .C2(n15528), .ZN(n25867) );
  NR4D0 U8664 ( .A1(n25871), .A2(n25872), .A3(n25873), .A4(n25874), .ZN(n25860) );
  OAI22D0 U8665 ( .A1(n24928), .A2(n3206), .B1(n24926), .B2(n3110), .ZN(n25874) );
  OAI222D0 U8666 ( .A1(n25002), .A2(n3446), .B1(n24929), .B2(n3254), .C1(
        n24933), .C2(n2342), .ZN(n25873) );
  OAI222D0 U8667 ( .A1(n25003), .A2(n3590), .B1(n25004), .B2(n3494), .C1(
        n25005), .C2(n3542), .ZN(n25872) );
  OAI222D0 U8668 ( .A1(n24965), .A2(n2582), .B1(n25006), .B2(n3638), .C1(
        n25007), .C2(n3686), .ZN(n25871) );
  NR4D0 U8669 ( .A1(n25875), .A2(n25876), .A3(n25877), .A4(n25878), .ZN(n25859) );
  OAI22D0 U8670 ( .A1(n25012), .A2(n5126), .B1(n24966), .B2(n2294), .ZN(n25878) );
  OAI222D0 U8671 ( .A1(n24925), .A2(n3062), .B1(n24923), .B2(n2966), .C1(
        n24960), .C2(n2870), .ZN(n25877) );
  OAI222D0 U8672 ( .A1(n25013), .A2(n5510), .B1(n25014), .B2(n5558), .C1(
        n24924), .C2(n3014), .ZN(n25876) );
  OAI222D0 U8673 ( .A1(n25015), .A2(n6086), .B1(n25016), .B2(n5990), .C1(
        n25017), .C2(n6134), .ZN(n25875) );
  INR4D0 U8674 ( .A1(n25879), .B1(n25880), .B2(n25881), .B3(n25882), .ZN(
        n25857) );
  OAI222D0 U8675 ( .A1(n25022), .A2(n5462), .B1(n25023), .B2(n6326), .C1(
        n25024), .C2(n5414), .ZN(n25882) );
  OAI222D0 U8676 ( .A1(n25025), .A2(n4502), .B1(n25026), .B2(n24619), .C1(
        n25027), .C2(n5606), .ZN(n25881) );
  OR4D0 U8677 ( .A1(n25883), .A2(n25884), .A3(n25885), .A4(n25886), .Z(n25880)
         );
  OAI222D0 U8678 ( .A1(n25032), .A2(n4598), .B1(n25033), .B2(n5318), .C1(
        n25034), .C2(n6230), .ZN(n25886) );
  OAI222D0 U8679 ( .A1(n25035), .A2(n6182), .B1(n25036), .B2(n4550), .C1(
        n25037), .C2(n5366), .ZN(n25885) );
  OAI22D0 U8680 ( .A1(n27119), .A2(n25038), .B1(n27118), .B2(n25039), .ZN(
        n25884) );
  OAI222D0 U8681 ( .A1(n24874), .A2(n25040), .B1(n25041), .B2(n5846), .C1(
        n25042), .C2(n5798), .ZN(n25883) );
  CKND0 U8682 ( .I(\Mem[44][20] ), .ZN(n24874) );
  AOI221D0 U8683 ( .A1(n27116), .A2(n25043), .B1(n27117), .B2(n25044), .C(
        n25887), .ZN(n25879) );
  OAI222D0 U8684 ( .A1(n25046), .A2(n6038), .B1(n24875), .B2(n25047), .C1(
        n25048), .C2(n4694), .ZN(n25887) );
  CKND0 U8685 ( .I(\Mem[45][20] ), .ZN(n24875) );
  NR4D0 U8686 ( .A1(n25888), .A2(n25889), .A3(n25890), .A4(n25891), .ZN(n25856) );
  OAI22D0 U8687 ( .A1(n25053), .A2(n5894), .B1(n25054), .B2(n5702), .ZN(n25891) );
  OAI222D0 U8688 ( .A1(n25055), .A2(n3830), .B1(n25056), .B2(n3878), .C1(
        n25057), .C2(n5942), .ZN(n25890) );
  OAI222D0 U8689 ( .A1(n25058), .A2(n3974), .B1(n25059), .B2(n4022), .C1(
        n25060), .C2(n3926), .ZN(n25889) );
  OAI222D0 U8690 ( .A1(n25061), .A2(n4118), .B1(n25062), .B2(n4166), .C1(
        n25063), .C2(n4070), .ZN(n25888) );
  NR4D0 U8691 ( .A1(n25892), .A2(n25893), .A3(n25894), .A4(n25895), .ZN(n25855) );
  OAI22D0 U8692 ( .A1(n25068), .A2(n2390), .B1(n25069), .B2(n2918), .ZN(n25895) );
  OAI222D0 U8693 ( .A1(n25070), .A2(n2486), .B1(n25071), .B2(n4310), .C1(
        n25072), .C2(n2630), .ZN(n25894) );
  OAI222D0 U8694 ( .A1(n25073), .A2(n4262), .B1(n24930), .B2(n3302), .C1(
        n25074), .C2(n4214), .ZN(n25893) );
  OAI222D0 U8695 ( .A1(n24932), .A2(n3398), .B1(n25075), .B2(n4838), .C1(
        n24931), .C2(n3350), .ZN(n25892) );
  ND4D0 U8696 ( .A1(n25896), .A2(n25897), .A3(n25898), .A4(n25899), .ZN(n2196)
         );
  AN4D0 U8697 ( .A1(n25900), .A2(n25901), .A3(n25902), .A4(n25903), .Z(n25899)
         );
  NR4D0 U8698 ( .A1(n25904), .A2(n25905), .A3(n25906), .A4(n25907), .ZN(n25903) );
  OAI222D0 U8699 ( .A1(n24979), .A2(n15533), .B1(n24980), .B2(n4453), .C1(
        n24964), .C2(n2245), .ZN(n25907) );
  OAI222D0 U8700 ( .A1(n24920), .A2(n2533), .B1(n24981), .B2(n5173), .C1(
        n24963), .C2(n2437), .ZN(n25906) );
  OAI222D0 U8701 ( .A1(n24982), .A2(n4933), .B1(n24983), .B2(n4981), .C1(
        n24984), .C2(n4885), .ZN(n25905) );
  OAI222D0 U8702 ( .A1(n24985), .A2(n4405), .B1(n24986), .B2(n3781), .C1(
        n24987), .C2(n4357), .ZN(n25904) );
  NR4D0 U8703 ( .A1(n25908), .A2(n25909), .A3(n25910), .A4(n25911), .ZN(n25902) );
  OAI22D0 U8704 ( .A1(n24922), .A2(n2821), .B1(n24992), .B2(n3733), .ZN(n25911) );
  OAI222D0 U8705 ( .A1(n24993), .A2(n17989), .B1(n24962), .B2(n2773), .C1(
        n24994), .C2(n17990), .ZN(n25910) );
  OAI222D0 U8706 ( .A1(n24995), .A2(n5221), .B1(n24961), .B2(n2677), .C1(
        n24921), .C2(n2725), .ZN(n25909) );
  OAI222D0 U8707 ( .A1(n24927), .A2(n3157), .B1(n24996), .B2(n4789), .C1(
        n24997), .C2(n15532), .ZN(n25908) );
  NR4D0 U8708 ( .A1(n25912), .A2(n25913), .A3(n25914), .A4(n25915), .ZN(n25901) );
  OAI22D0 U8709 ( .A1(n24928), .A2(n3205), .B1(n24926), .B2(n3109), .ZN(n25915) );
  OAI222D0 U8710 ( .A1(n25002), .A2(n3445), .B1(n24929), .B2(n3253), .C1(
        n24933), .C2(n2341), .ZN(n25914) );
  OAI222D0 U8711 ( .A1(n25003), .A2(n3589), .B1(n25004), .B2(n3493), .C1(
        n25005), .C2(n3541), .ZN(n25913) );
  OAI222D0 U8712 ( .A1(n24965), .A2(n2581), .B1(n25006), .B2(n3637), .C1(
        n25007), .C2(n3685), .ZN(n25912) );
  NR4D0 U8713 ( .A1(n25916), .A2(n25917), .A3(n25918), .A4(n25919), .ZN(n25900) );
  OAI22D0 U8714 ( .A1(n25012), .A2(n5125), .B1(n24966), .B2(n2293), .ZN(n25919) );
  OAI222D0 U8715 ( .A1(n24925), .A2(n3061), .B1(n24923), .B2(n2965), .C1(
        n24960), .C2(n2869), .ZN(n25918) );
  OAI222D0 U8716 ( .A1(n25013), .A2(n5509), .B1(n25014), .B2(n5557), .C1(
        n24924), .C2(n3013), .ZN(n25917) );
  OAI222D0 U8717 ( .A1(n25015), .A2(n6085), .B1(n25016), .B2(n5989), .C1(
        n25017), .C2(n6133), .ZN(n25916) );
  INR4D0 U8718 ( .A1(n25920), .B1(n25921), .B2(n25922), .B3(n25923), .ZN(
        n25898) );
  OAI222D0 U8719 ( .A1(n25022), .A2(n5461), .B1(n25023), .B2(n6325), .C1(
        n25024), .C2(n5413), .ZN(n25923) );
  OAI222D0 U8720 ( .A1(n25025), .A2(n4501), .B1(n25026), .B2(n24622), .C1(
        n25027), .C2(n5605), .ZN(n25922) );
  OR4D0 U8721 ( .A1(n25924), .A2(n25925), .A3(n25926), .A4(n25927), .Z(n25921)
         );
  OAI222D0 U8722 ( .A1(n25032), .A2(n4597), .B1(n25033), .B2(n5317), .C1(
        n25034), .C2(n6229), .ZN(n25927) );
  OAI222D0 U8723 ( .A1(n25035), .A2(n6181), .B1(n25036), .B2(n4549), .C1(
        n25037), .C2(n5365), .ZN(n25926) );
  OAI22D0 U8724 ( .A1(n27123), .A2(n25038), .B1(n27122), .B2(n25039), .ZN(
        n25925) );
  OAI222D0 U8725 ( .A1(n24872), .A2(n25040), .B1(n25041), .B2(n5845), .C1(
        n25042), .C2(n5797), .ZN(n25924) );
  CKND0 U8726 ( .I(\Mem[44][21] ), .ZN(n24872) );
  AOI221D0 U8727 ( .A1(n27120), .A2(n25043), .B1(n27121), .B2(n25044), .C(
        n25928), .ZN(n25920) );
  OAI222D0 U8728 ( .A1(n25046), .A2(n6037), .B1(n24873), .B2(n25047), .C1(
        n25048), .C2(n4693), .ZN(n25928) );
  CKND0 U8729 ( .I(\Mem[45][21] ), .ZN(n24873) );
  NR4D0 U8730 ( .A1(n25929), .A2(n25930), .A3(n25931), .A4(n25932), .ZN(n25897) );
  OAI22D0 U8731 ( .A1(n25053), .A2(n5893), .B1(n25054), .B2(n5701), .ZN(n25932) );
  OAI222D0 U8732 ( .A1(n25055), .A2(n3829), .B1(n25056), .B2(n3877), .C1(
        n25057), .C2(n5941), .ZN(n25931) );
  OAI222D0 U8733 ( .A1(n25058), .A2(n3973), .B1(n25059), .B2(n4021), .C1(
        n25060), .C2(n3925), .ZN(n25930) );
  OAI222D0 U8734 ( .A1(n25061), .A2(n4117), .B1(n25062), .B2(n4165), .C1(
        n25063), .C2(n4069), .ZN(n25929) );
  NR4D0 U8735 ( .A1(n25933), .A2(n25934), .A3(n25935), .A4(n25936), .ZN(n25896) );
  OAI22D0 U8736 ( .A1(n25068), .A2(n2389), .B1(n25069), .B2(n2917), .ZN(n25936) );
  OAI222D0 U8737 ( .A1(n25070), .A2(n2485), .B1(n25071), .B2(n4309), .C1(
        n25072), .C2(n2629), .ZN(n25935) );
  OAI222D0 U8738 ( .A1(n25073), .A2(n4261), .B1(n24930), .B2(n3301), .C1(
        n25074), .C2(n4213), .ZN(n25934) );
  OAI222D0 U8739 ( .A1(n24932), .A2(n3397), .B1(n25075), .B2(n4837), .C1(
        n24931), .C2(n3349), .ZN(n25933) );
  ND4D0 U8740 ( .A1(n25937), .A2(n25938), .A3(n25939), .A4(n25940), .ZN(n2195)
         );
  AN4D0 U8741 ( .A1(n25941), .A2(n25942), .A3(n25943), .A4(n25944), .Z(n25940)
         );
  NR4D0 U8742 ( .A1(n25945), .A2(n25946), .A3(n25947), .A4(n25948), .ZN(n25944) );
  OAI222D0 U8743 ( .A1(n24979), .A2(n15537), .B1(n24980), .B2(n4452), .C1(
        n24964), .C2(n2244), .ZN(n25948) );
  OAI222D0 U8744 ( .A1(n24920), .A2(n2532), .B1(n24981), .B2(n5172), .C1(
        n24963), .C2(n2436), .ZN(n25947) );
  OAI222D0 U8745 ( .A1(n24982), .A2(n4932), .B1(n24983), .B2(n4980), .C1(
        n24984), .C2(n4884), .ZN(n25946) );
  OAI222D0 U8746 ( .A1(n24985), .A2(n4404), .B1(n24986), .B2(n3780), .C1(
        n24987), .C2(n4356), .ZN(n25945) );
  NR4D0 U8747 ( .A1(n25949), .A2(n25950), .A3(n25951), .A4(n25952), .ZN(n25943) );
  OAI22D0 U8748 ( .A1(n24922), .A2(n2820), .B1(n24992), .B2(n3732), .ZN(n25952) );
  OAI222D0 U8749 ( .A1(n24993), .A2(n17992), .B1(n24962), .B2(n2772), .C1(
        n24994), .C2(n17993), .ZN(n25951) );
  OAI222D0 U8750 ( .A1(n24995), .A2(n5220), .B1(n24961), .B2(n2676), .C1(
        n24921), .C2(n2724), .ZN(n25950) );
  OAI222D0 U8751 ( .A1(n24927), .A2(n3156), .B1(n24996), .B2(n4788), .C1(
        n24997), .C2(n15536), .ZN(n25949) );
  NR4D0 U8752 ( .A1(n25953), .A2(n25954), .A3(n25955), .A4(n25956), .ZN(n25942) );
  OAI22D0 U8753 ( .A1(n24928), .A2(n3204), .B1(n24926), .B2(n3108), .ZN(n25956) );
  OAI222D0 U8754 ( .A1(n25002), .A2(n3444), .B1(n24929), .B2(n3252), .C1(
        n24933), .C2(n2340), .ZN(n25955) );
  OAI222D0 U8755 ( .A1(n25003), .A2(n3588), .B1(n25004), .B2(n3492), .C1(
        n25005), .C2(n3540), .ZN(n25954) );
  OAI222D0 U8756 ( .A1(n24965), .A2(n2580), .B1(n25006), .B2(n3636), .C1(
        n25007), .C2(n3684), .ZN(n25953) );
  NR4D0 U8757 ( .A1(n25957), .A2(n25958), .A3(n25959), .A4(n25960), .ZN(n25941) );
  OAI22D0 U8758 ( .A1(n25012), .A2(n5124), .B1(n24966), .B2(n2292), .ZN(n25960) );
  OAI222D0 U8759 ( .A1(n24925), .A2(n3060), .B1(n24923), .B2(n2964), .C1(
        n24960), .C2(n2868), .ZN(n25959) );
  OAI222D0 U8760 ( .A1(n25013), .A2(n5508), .B1(n25014), .B2(n5556), .C1(
        n24924), .C2(n3012), .ZN(n25958) );
  OAI222D0 U8761 ( .A1(n25015), .A2(n6084), .B1(n25016), .B2(n5988), .C1(
        n25017), .C2(n6132), .ZN(n25957) );
  INR4D0 U8762 ( .A1(n25961), .B1(n25962), .B2(n25963), .B3(n25964), .ZN(
        n25939) );
  OAI222D0 U8763 ( .A1(n25022), .A2(n5460), .B1(n25023), .B2(n6324), .C1(
        n25024), .C2(n5412), .ZN(n25964) );
  OAI222D0 U8764 ( .A1(n25025), .A2(n4500), .B1(n25026), .B2(n24625), .C1(
        n25027), .C2(n5604), .ZN(n25963) );
  OR4D0 U8765 ( .A1(n25965), .A2(n25966), .A3(n25967), .A4(n25968), .Z(n25962)
         );
  OAI222D0 U8766 ( .A1(n25032), .A2(n4596), .B1(n25033), .B2(n5316), .C1(
        n25034), .C2(n6228), .ZN(n25968) );
  OAI222D0 U8767 ( .A1(n25035), .A2(n6180), .B1(n25036), .B2(n4548), .C1(
        n25037), .C2(n5364), .ZN(n25967) );
  OAI22D0 U8768 ( .A1(n27127), .A2(n25038), .B1(n27126), .B2(n25039), .ZN(
        n25966) );
  OAI222D0 U8769 ( .A1(n24870), .A2(n25040), .B1(n25041), .B2(n5844), .C1(
        n25042), .C2(n5796), .ZN(n25965) );
  CKND0 U8770 ( .I(\Mem[44][22] ), .ZN(n24870) );
  AOI221D0 U8771 ( .A1(n27124), .A2(n25043), .B1(n27125), .B2(n25044), .C(
        n25969), .ZN(n25961) );
  OAI222D0 U8772 ( .A1(n25046), .A2(n6036), .B1(n24871), .B2(n25047), .C1(
        n25048), .C2(n4692), .ZN(n25969) );
  CKND0 U8773 ( .I(\Mem[45][22] ), .ZN(n24871) );
  NR4D0 U8774 ( .A1(n25970), .A2(n25971), .A3(n25972), .A4(n25973), .ZN(n25938) );
  OAI22D0 U8775 ( .A1(n25053), .A2(n5892), .B1(n25054), .B2(n5700), .ZN(n25973) );
  OAI222D0 U8776 ( .A1(n25055), .A2(n3828), .B1(n25056), .B2(n3876), .C1(
        n25057), .C2(n5940), .ZN(n25972) );
  OAI222D0 U8777 ( .A1(n25058), .A2(n3972), .B1(n25059), .B2(n4020), .C1(
        n25060), .C2(n3924), .ZN(n25971) );
  OAI222D0 U8778 ( .A1(n25061), .A2(n4116), .B1(n25062), .B2(n4164), .C1(
        n25063), .C2(n4068), .ZN(n25970) );
  NR4D0 U8779 ( .A1(n25974), .A2(n25975), .A3(n25976), .A4(n25977), .ZN(n25937) );
  OAI22D0 U8780 ( .A1(n25068), .A2(n2388), .B1(n25069), .B2(n2916), .ZN(n25977) );
  OAI222D0 U8781 ( .A1(n25070), .A2(n2484), .B1(n25071), .B2(n4308), .C1(
        n25072), .C2(n2628), .ZN(n25976) );
  OAI222D0 U8782 ( .A1(n25073), .A2(n4260), .B1(n24930), .B2(n3300), .C1(
        n25074), .C2(n4212), .ZN(n25975) );
  OAI222D0 U8783 ( .A1(n24932), .A2(n3396), .B1(n25075), .B2(n4836), .C1(
        n24931), .C2(n3348), .ZN(n25974) );
  ND4D0 U8784 ( .A1(n25978), .A2(n25979), .A3(n25980), .A4(n25981), .ZN(n2194)
         );
  AN4D0 U8785 ( .A1(n25982), .A2(n25983), .A3(n25984), .A4(n25985), .Z(n25981)
         );
  NR4D0 U8786 ( .A1(n25986), .A2(n25987), .A3(n25988), .A4(n25989), .ZN(n25985) );
  OAI222D0 U8787 ( .A1(n24979), .A2(n15541), .B1(n24980), .B2(n4451), .C1(
        n24964), .C2(n2243), .ZN(n25989) );
  OAI222D0 U8788 ( .A1(n24920), .A2(n2531), .B1(n24981), .B2(n5171), .C1(
        n24963), .C2(n2435), .ZN(n25988) );
  OAI222D0 U8789 ( .A1(n24982), .A2(n4931), .B1(n24983), .B2(n4979), .C1(
        n24984), .C2(n4883), .ZN(n25987) );
  OAI222D0 U8790 ( .A1(n24985), .A2(n4403), .B1(n24986), .B2(n3779), .C1(
        n24987), .C2(n4355), .ZN(n25986) );
  NR4D0 U8791 ( .A1(n25990), .A2(n25991), .A3(n25992), .A4(n25993), .ZN(n25984) );
  OAI22D0 U8792 ( .A1(n24922), .A2(n2819), .B1(n24992), .B2(n3731), .ZN(n25993) );
  OAI222D0 U8793 ( .A1(n24993), .A2(n17995), .B1(n24962), .B2(n2771), .C1(
        n24994), .C2(n17996), .ZN(n25992) );
  OAI222D0 U8794 ( .A1(n24995), .A2(n5219), .B1(n24961), .B2(n2675), .C1(
        n24921), .C2(n2723), .ZN(n25991) );
  OAI222D0 U8795 ( .A1(n24927), .A2(n3155), .B1(n24996), .B2(n4787), .C1(
        n24997), .C2(n15540), .ZN(n25990) );
  NR4D0 U8796 ( .A1(n25994), .A2(n25995), .A3(n25996), .A4(n25997), .ZN(n25983) );
  OAI22D0 U8797 ( .A1(n24928), .A2(n3203), .B1(n24926), .B2(n3107), .ZN(n25997) );
  OAI222D0 U8798 ( .A1(n25002), .A2(n3443), .B1(n24929), .B2(n3251), .C1(
        n24933), .C2(n2339), .ZN(n25996) );
  OAI222D0 U8799 ( .A1(n25003), .A2(n3587), .B1(n25004), .B2(n3491), .C1(
        n25005), .C2(n3539), .ZN(n25995) );
  OAI222D0 U8800 ( .A1(n24965), .A2(n2579), .B1(n25006), .B2(n3635), .C1(
        n25007), .C2(n3683), .ZN(n25994) );
  NR4D0 U8801 ( .A1(n25998), .A2(n25999), .A3(n26000), .A4(n26001), .ZN(n25982) );
  OAI22D0 U8802 ( .A1(n25012), .A2(n5123), .B1(n24966), .B2(n2291), .ZN(n26001) );
  OAI222D0 U8803 ( .A1(n24925), .A2(n3059), .B1(n24923), .B2(n2963), .C1(
        n24960), .C2(n2867), .ZN(n26000) );
  OAI222D0 U8804 ( .A1(n25013), .A2(n5507), .B1(n25014), .B2(n5555), .C1(
        n24924), .C2(n3011), .ZN(n25999) );
  OAI222D0 U8805 ( .A1(n25015), .A2(n6083), .B1(n25016), .B2(n5987), .C1(
        n25017), .C2(n6131), .ZN(n25998) );
  INR4D0 U8806 ( .A1(n26002), .B1(n26003), .B2(n26004), .B3(n26005), .ZN(
        n25980) );
  OAI222D0 U8807 ( .A1(n25022), .A2(n5459), .B1(n25023), .B2(n6323), .C1(
        n25024), .C2(n5411), .ZN(n26005) );
  OAI222D0 U8808 ( .A1(n25025), .A2(n4499), .B1(n25026), .B2(n24628), .C1(
        n25027), .C2(n5603), .ZN(n26004) );
  OR4D0 U8809 ( .A1(n26006), .A2(n26007), .A3(n26008), .A4(n26009), .Z(n26003)
         );
  OAI222D0 U8810 ( .A1(n25032), .A2(n4595), .B1(n25033), .B2(n5315), .C1(
        n25034), .C2(n6227), .ZN(n26009) );
  OAI222D0 U8811 ( .A1(n25035), .A2(n6179), .B1(n25036), .B2(n4547), .C1(
        n25037), .C2(n5363), .ZN(n26008) );
  OAI22D0 U8812 ( .A1(n27131), .A2(n25038), .B1(n27130), .B2(n25039), .ZN(
        n26007) );
  OAI222D0 U8813 ( .A1(n24868), .A2(n25040), .B1(n25041), .B2(n5843), .C1(
        n25042), .C2(n5795), .ZN(n26006) );
  CKND0 U8814 ( .I(\Mem[44][23] ), .ZN(n24868) );
  AOI221D0 U8815 ( .A1(n27128), .A2(n25043), .B1(n27129), .B2(n25044), .C(
        n26010), .ZN(n26002) );
  OAI222D0 U8816 ( .A1(n25046), .A2(n6035), .B1(n24869), .B2(n25047), .C1(
        n25048), .C2(n4691), .ZN(n26010) );
  CKND0 U8817 ( .I(\Mem[45][23] ), .ZN(n24869) );
  NR4D0 U8818 ( .A1(n26011), .A2(n26012), .A3(n26013), .A4(n26014), .ZN(n25979) );
  OAI22D0 U8819 ( .A1(n25053), .A2(n5891), .B1(n25054), .B2(n5699), .ZN(n26014) );
  OAI222D0 U8820 ( .A1(n25055), .A2(n3827), .B1(n25056), .B2(n3875), .C1(
        n25057), .C2(n5939), .ZN(n26013) );
  OAI222D0 U8821 ( .A1(n25058), .A2(n3971), .B1(n25059), .B2(n4019), .C1(
        n25060), .C2(n3923), .ZN(n26012) );
  OAI222D0 U8822 ( .A1(n25061), .A2(n4115), .B1(n25062), .B2(n4163), .C1(
        n25063), .C2(n4067), .ZN(n26011) );
  NR4D0 U8823 ( .A1(n26015), .A2(n26016), .A3(n26017), .A4(n26018), .ZN(n25978) );
  OAI22D0 U8824 ( .A1(n25068), .A2(n2387), .B1(n25069), .B2(n2915), .ZN(n26018) );
  OAI222D0 U8825 ( .A1(n25070), .A2(n2483), .B1(n25071), .B2(n4307), .C1(
        n25072), .C2(n2627), .ZN(n26017) );
  OAI222D0 U8826 ( .A1(n25073), .A2(n4259), .B1(n24930), .B2(n3299), .C1(
        n25074), .C2(n4211), .ZN(n26016) );
  OAI222D0 U8827 ( .A1(n24932), .A2(n3395), .B1(n25075), .B2(n4835), .C1(
        n24931), .C2(n3347), .ZN(n26015) );
  ND4D0 U8828 ( .A1(n26019), .A2(n26020), .A3(n26021), .A4(n26022), .ZN(n2193)
         );
  AN4D0 U8829 ( .A1(n26023), .A2(n26024), .A3(n26025), .A4(n26026), .Z(n26022)
         );
  NR4D0 U8830 ( .A1(n26027), .A2(n26028), .A3(n26029), .A4(n26030), .ZN(n26026) );
  OAI222D0 U8831 ( .A1(n24979), .A2(n15545), .B1(n24980), .B2(n4450), .C1(
        n24964), .C2(n2242), .ZN(n26030) );
  OAI222D0 U8832 ( .A1(n24920), .A2(n2530), .B1(n24981), .B2(n5170), .C1(
        n24963), .C2(n2434), .ZN(n26029) );
  OAI222D0 U8833 ( .A1(n24982), .A2(n4930), .B1(n24983), .B2(n4978), .C1(
        n24984), .C2(n4882), .ZN(n26028) );
  OAI222D0 U8834 ( .A1(n24985), .A2(n4402), .B1(n24986), .B2(n3778), .C1(
        n24987), .C2(n4354), .ZN(n26027) );
  NR4D0 U8835 ( .A1(n26031), .A2(n26032), .A3(n26033), .A4(n26034), .ZN(n26025) );
  OAI22D0 U8836 ( .A1(n24922), .A2(n2818), .B1(n24992), .B2(n3730), .ZN(n26034) );
  OAI222D0 U8837 ( .A1(n24993), .A2(n17998), .B1(n24962), .B2(n2770), .C1(
        n24994), .C2(n17999), .ZN(n26033) );
  OAI222D0 U8838 ( .A1(n24995), .A2(n5218), .B1(n24961), .B2(n2674), .C1(
        n24921), .C2(n2722), .ZN(n26032) );
  OAI222D0 U8839 ( .A1(n24927), .A2(n3154), .B1(n24996), .B2(n4786), .C1(
        n24997), .C2(n15544), .ZN(n26031) );
  NR4D0 U8840 ( .A1(n26035), .A2(n26036), .A3(n26037), .A4(n26038), .ZN(n26024) );
  OAI22D0 U8841 ( .A1(n24928), .A2(n3202), .B1(n24926), .B2(n3106), .ZN(n26038) );
  OAI222D0 U8842 ( .A1(n25002), .A2(n3442), .B1(n24929), .B2(n3250), .C1(
        n24933), .C2(n2338), .ZN(n26037) );
  OAI222D0 U8843 ( .A1(n25003), .A2(n3586), .B1(n25004), .B2(n3490), .C1(
        n25005), .C2(n3538), .ZN(n26036) );
  OAI222D0 U8844 ( .A1(n24965), .A2(n2578), .B1(n25006), .B2(n3634), .C1(
        n25007), .C2(n3682), .ZN(n26035) );
  NR4D0 U8845 ( .A1(n26039), .A2(n26040), .A3(n26041), .A4(n26042), .ZN(n26023) );
  OAI22D0 U8846 ( .A1(n25012), .A2(n5122), .B1(n24966), .B2(n2290), .ZN(n26042) );
  OAI222D0 U8847 ( .A1(n24925), .A2(n3058), .B1(n24923), .B2(n2962), .C1(
        n24960), .C2(n2866), .ZN(n26041) );
  OAI222D0 U8848 ( .A1(n25013), .A2(n5506), .B1(n25014), .B2(n5554), .C1(
        n24924), .C2(n3010), .ZN(n26040) );
  OAI222D0 U8849 ( .A1(n25015), .A2(n6082), .B1(n25016), .B2(n5986), .C1(
        n25017), .C2(n6130), .ZN(n26039) );
  INR4D0 U8850 ( .A1(n26043), .B1(n26044), .B2(n26045), .B3(n26046), .ZN(
        n26021) );
  OAI222D0 U8851 ( .A1(n25022), .A2(n5458), .B1(n25023), .B2(n6322), .C1(
        n25024), .C2(n5410), .ZN(n26046) );
  OAI222D0 U8852 ( .A1(n25025), .A2(n4498), .B1(n25026), .B2(n24631), .C1(
        n25027), .C2(n5602), .ZN(n26045) );
  OR4D0 U8853 ( .A1(n26047), .A2(n26048), .A3(n26049), .A4(n26050), .Z(n26044)
         );
  OAI222D0 U8854 ( .A1(n25032), .A2(n4594), .B1(n25033), .B2(n5314), .C1(
        n25034), .C2(n6226), .ZN(n26050) );
  OAI222D0 U8855 ( .A1(n25035), .A2(n6178), .B1(n25036), .B2(n4546), .C1(
        n25037), .C2(n5362), .ZN(n26049) );
  OAI22D0 U8856 ( .A1(n27135), .A2(n25038), .B1(n27134), .B2(n25039), .ZN(
        n26048) );
  OAI222D0 U8857 ( .A1(n24866), .A2(n25040), .B1(n25041), .B2(n5842), .C1(
        n25042), .C2(n5794), .ZN(n26047) );
  CKND0 U8858 ( .I(\Mem[44][24] ), .ZN(n24866) );
  AOI221D0 U8859 ( .A1(n27132), .A2(n25043), .B1(n27133), .B2(n25044), .C(
        n26051), .ZN(n26043) );
  OAI222D0 U8860 ( .A1(n25046), .A2(n6034), .B1(n24867), .B2(n25047), .C1(
        n25048), .C2(n4690), .ZN(n26051) );
  CKND0 U8861 ( .I(\Mem[45][24] ), .ZN(n24867) );
  NR4D0 U8862 ( .A1(n26052), .A2(n26053), .A3(n26054), .A4(n26055), .ZN(n26020) );
  OAI22D0 U8863 ( .A1(n25053), .A2(n5890), .B1(n25054), .B2(n5698), .ZN(n26055) );
  OAI222D0 U8864 ( .A1(n25055), .A2(n3826), .B1(n25056), .B2(n3874), .C1(
        n25057), .C2(n5938), .ZN(n26054) );
  OAI222D0 U8865 ( .A1(n25058), .A2(n3970), .B1(n25059), .B2(n4018), .C1(
        n25060), .C2(n3922), .ZN(n26053) );
  OAI222D0 U8866 ( .A1(n25061), .A2(n4114), .B1(n25062), .B2(n4162), .C1(
        n25063), .C2(n4066), .ZN(n26052) );
  NR4D0 U8867 ( .A1(n26056), .A2(n26057), .A3(n26058), .A4(n26059), .ZN(n26019) );
  OAI22D0 U8868 ( .A1(n25068), .A2(n2386), .B1(n25069), .B2(n2914), .ZN(n26059) );
  OAI222D0 U8869 ( .A1(n25070), .A2(n2482), .B1(n25071), .B2(n4306), .C1(
        n25072), .C2(n2626), .ZN(n26058) );
  OAI222D0 U8870 ( .A1(n25073), .A2(n4258), .B1(n24930), .B2(n3298), .C1(
        n25074), .C2(n4210), .ZN(n26057) );
  OAI222D0 U8871 ( .A1(n24932), .A2(n3394), .B1(n25075), .B2(n4834), .C1(
        n24931), .C2(n3346), .ZN(n26056) );
  ND4D0 U8872 ( .A1(n26060), .A2(n26061), .A3(n26062), .A4(n26063), .ZN(n2192)
         );
  AN4D0 U8873 ( .A1(n26064), .A2(n26065), .A3(n26066), .A4(n26067), .Z(n26063)
         );
  NR4D0 U8874 ( .A1(n26068), .A2(n26069), .A3(n26070), .A4(n26071), .ZN(n26067) );
  OAI222D0 U8875 ( .A1(n24979), .A2(n15549), .B1(n24980), .B2(n4449), .C1(
        n24964), .C2(n2241), .ZN(n26071) );
  OAI222D0 U8876 ( .A1(n24920), .A2(n2529), .B1(n24981), .B2(n5169), .C1(
        n24963), .C2(n2433), .ZN(n26070) );
  OAI222D0 U8877 ( .A1(n24982), .A2(n4929), .B1(n24983), .B2(n4977), .C1(
        n24984), .C2(n4881), .ZN(n26069) );
  OAI222D0 U8878 ( .A1(n24985), .A2(n4401), .B1(n24986), .B2(n3777), .C1(
        n24987), .C2(n4353), .ZN(n26068) );
  NR4D0 U8879 ( .A1(n26072), .A2(n26073), .A3(n26074), .A4(n26075), .ZN(n26066) );
  OAI22D0 U8880 ( .A1(n24922), .A2(n2817), .B1(n24992), .B2(n3729), .ZN(n26075) );
  OAI222D0 U8881 ( .A1(n24993), .A2(n18001), .B1(n24962), .B2(n2769), .C1(
        n24994), .C2(n18002), .ZN(n26074) );
  OAI222D0 U8882 ( .A1(n24995), .A2(n5217), .B1(n24961), .B2(n2673), .C1(
        n24921), .C2(n2721), .ZN(n26073) );
  OAI222D0 U8883 ( .A1(n24927), .A2(n3153), .B1(n24996), .B2(n4785), .C1(
        n24997), .C2(n15548), .ZN(n26072) );
  NR4D0 U8884 ( .A1(n26076), .A2(n26077), .A3(n26078), .A4(n26079), .ZN(n26065) );
  OAI22D0 U8885 ( .A1(n24928), .A2(n3201), .B1(n24926), .B2(n3105), .ZN(n26079) );
  OAI222D0 U8886 ( .A1(n25002), .A2(n3441), .B1(n24929), .B2(n3249), .C1(
        n24933), .C2(n2337), .ZN(n26078) );
  OAI222D0 U8887 ( .A1(n25003), .A2(n3585), .B1(n25004), .B2(n3489), .C1(
        n25005), .C2(n3537), .ZN(n26077) );
  OAI222D0 U8888 ( .A1(n24965), .A2(n2577), .B1(n25006), .B2(n3633), .C1(
        n25007), .C2(n3681), .ZN(n26076) );
  NR4D0 U8889 ( .A1(n26080), .A2(n26081), .A3(n26082), .A4(n26083), .ZN(n26064) );
  OAI22D0 U8890 ( .A1(n25012), .A2(n5121), .B1(n24966), .B2(n2289), .ZN(n26083) );
  OAI222D0 U8891 ( .A1(n24925), .A2(n3057), .B1(n24923), .B2(n2961), .C1(
        n24960), .C2(n2865), .ZN(n26082) );
  OAI222D0 U8892 ( .A1(n25013), .A2(n5505), .B1(n25014), .B2(n5553), .C1(
        n24924), .C2(n3009), .ZN(n26081) );
  OAI222D0 U8893 ( .A1(n25015), .A2(n6081), .B1(n25016), .B2(n5985), .C1(
        n25017), .C2(n6129), .ZN(n26080) );
  INR4D0 U8894 ( .A1(n26084), .B1(n26085), .B2(n26086), .B3(n26087), .ZN(
        n26062) );
  OAI222D0 U8895 ( .A1(n25022), .A2(n5457), .B1(n25023), .B2(n6321), .C1(
        n25024), .C2(n5409), .ZN(n26087) );
  OAI222D0 U8896 ( .A1(n25025), .A2(n4497), .B1(n25026), .B2(n24634), .C1(
        n25027), .C2(n5601), .ZN(n26086) );
  OR4D0 U8897 ( .A1(n26088), .A2(n26089), .A3(n26090), .A4(n26091), .Z(n26085)
         );
  OAI222D0 U8898 ( .A1(n25032), .A2(n4593), .B1(n25033), .B2(n5313), .C1(
        n25034), .C2(n6225), .ZN(n26091) );
  OAI222D0 U8899 ( .A1(n25035), .A2(n6177), .B1(n25036), .B2(n4545), .C1(
        n25037), .C2(n5361), .ZN(n26090) );
  OAI22D0 U8900 ( .A1(n27139), .A2(n25038), .B1(n27138), .B2(n25039), .ZN(
        n26089) );
  OAI222D0 U8901 ( .A1(n24864), .A2(n25040), .B1(n25041), .B2(n5841), .C1(
        n25042), .C2(n5793), .ZN(n26088) );
  CKND0 U8902 ( .I(\Mem[44][25] ), .ZN(n24864) );
  AOI221D0 U8903 ( .A1(n27136), .A2(n25043), .B1(n27137), .B2(n25044), .C(
        n26092), .ZN(n26084) );
  OAI222D0 U8904 ( .A1(n25046), .A2(n6033), .B1(n24865), .B2(n25047), .C1(
        n25048), .C2(n4689), .ZN(n26092) );
  CKND0 U8905 ( .I(\Mem[45][25] ), .ZN(n24865) );
  NR4D0 U8906 ( .A1(n26093), .A2(n26094), .A3(n26095), .A4(n26096), .ZN(n26061) );
  OAI22D0 U8907 ( .A1(n25053), .A2(n5889), .B1(n25054), .B2(n5697), .ZN(n26096) );
  OAI222D0 U8908 ( .A1(n25055), .A2(n3825), .B1(n25056), .B2(n3873), .C1(
        n25057), .C2(n5937), .ZN(n26095) );
  OAI222D0 U8909 ( .A1(n25058), .A2(n3969), .B1(n25059), .B2(n4017), .C1(
        n25060), .C2(n3921), .ZN(n26094) );
  OAI222D0 U8910 ( .A1(n25061), .A2(n4113), .B1(n25062), .B2(n4161), .C1(
        n25063), .C2(n4065), .ZN(n26093) );
  NR4D0 U8911 ( .A1(n26097), .A2(n26098), .A3(n26099), .A4(n26100), .ZN(n26060) );
  OAI22D0 U8912 ( .A1(n25068), .A2(n2385), .B1(n25069), .B2(n2913), .ZN(n26100) );
  OAI222D0 U8913 ( .A1(n25070), .A2(n2481), .B1(n25071), .B2(n4305), .C1(
        n25072), .C2(n2625), .ZN(n26099) );
  OAI222D0 U8914 ( .A1(n25073), .A2(n4257), .B1(n24930), .B2(n3297), .C1(
        n25074), .C2(n4209), .ZN(n26098) );
  OAI222D0 U8915 ( .A1(n24932), .A2(n3393), .B1(n25075), .B2(n4833), .C1(
        n24931), .C2(n3345), .ZN(n26097) );
  ND4D0 U8916 ( .A1(n26101), .A2(n26102), .A3(n26103), .A4(n26104), .ZN(n2191)
         );
  AN4D0 U8917 ( .A1(n26105), .A2(n26106), .A3(n26107), .A4(n26108), .Z(n26104)
         );
  NR4D0 U8918 ( .A1(n26109), .A2(n26110), .A3(n26111), .A4(n26112), .ZN(n26108) );
  OAI222D0 U8919 ( .A1(n24979), .A2(n15553), .B1(n24980), .B2(n4448), .C1(
        n24964), .C2(n2240), .ZN(n26112) );
  OAI222D0 U8920 ( .A1(n24920), .A2(n2528), .B1(n24981), .B2(n5168), .C1(
        n24963), .C2(n2432), .ZN(n26111) );
  OAI222D0 U8921 ( .A1(n24982), .A2(n4928), .B1(n24983), .B2(n4976), .C1(
        n24984), .C2(n4880), .ZN(n26110) );
  OAI222D0 U8922 ( .A1(n24985), .A2(n4400), .B1(n24986), .B2(n3776), .C1(
        n24987), .C2(n4352), .ZN(n26109) );
  NR4D0 U8923 ( .A1(n26113), .A2(n26114), .A3(n26115), .A4(n26116), .ZN(n26107) );
  OAI22D0 U8924 ( .A1(n24922), .A2(n2816), .B1(n24992), .B2(n3728), .ZN(n26116) );
  OAI222D0 U8925 ( .A1(n24993), .A2(n18004), .B1(n24962), .B2(n2768), .C1(
        n24994), .C2(n18005), .ZN(n26115) );
  OAI222D0 U8926 ( .A1(n24995), .A2(n5216), .B1(n24961), .B2(n2672), .C1(
        n24921), .C2(n2720), .ZN(n26114) );
  OAI222D0 U8927 ( .A1(n24927), .A2(n3152), .B1(n24996), .B2(n4784), .C1(
        n24997), .C2(n15552), .ZN(n26113) );
  NR4D0 U8928 ( .A1(n26117), .A2(n26118), .A3(n26119), .A4(n26120), .ZN(n26106) );
  OAI22D0 U8929 ( .A1(n24928), .A2(n3200), .B1(n24926), .B2(n3104), .ZN(n26120) );
  OAI222D0 U8930 ( .A1(n25002), .A2(n3440), .B1(n24929), .B2(n3248), .C1(
        n24933), .C2(n2336), .ZN(n26119) );
  OAI222D0 U8931 ( .A1(n25003), .A2(n3584), .B1(n25004), .B2(n3488), .C1(
        n25005), .C2(n3536), .ZN(n26118) );
  OAI222D0 U8932 ( .A1(n24965), .A2(n2576), .B1(n25006), .B2(n3632), .C1(
        n25007), .C2(n3680), .ZN(n26117) );
  NR4D0 U8933 ( .A1(n26121), .A2(n26122), .A3(n26123), .A4(n26124), .ZN(n26105) );
  OAI22D0 U8934 ( .A1(n25012), .A2(n5120), .B1(n24966), .B2(n2288), .ZN(n26124) );
  OAI222D0 U8935 ( .A1(n24925), .A2(n3056), .B1(n24923), .B2(n2960), .C1(
        n24960), .C2(n2864), .ZN(n26123) );
  OAI222D0 U8936 ( .A1(n25013), .A2(n5504), .B1(n25014), .B2(n5552), .C1(
        n24924), .C2(n3008), .ZN(n26122) );
  OAI222D0 U8937 ( .A1(n25015), .A2(n6080), .B1(n25016), .B2(n5984), .C1(
        n25017), .C2(n6128), .ZN(n26121) );
  INR4D0 U8938 ( .A1(n26125), .B1(n26126), .B2(n26127), .B3(n26128), .ZN(
        n26103) );
  OAI222D0 U8939 ( .A1(n25022), .A2(n5456), .B1(n25023), .B2(n6320), .C1(
        n25024), .C2(n5408), .ZN(n26128) );
  OAI222D0 U8940 ( .A1(n25025), .A2(n4496), .B1(n25026), .B2(n24637), .C1(
        n25027), .C2(n5600), .ZN(n26127) );
  OR4D0 U8941 ( .A1(n26129), .A2(n26130), .A3(n26131), .A4(n26132), .Z(n26126)
         );
  OAI222D0 U8942 ( .A1(n25032), .A2(n4592), .B1(n25033), .B2(n5312), .C1(
        n25034), .C2(n6224), .ZN(n26132) );
  OAI222D0 U8943 ( .A1(n25035), .A2(n6176), .B1(n25036), .B2(n4544), .C1(
        n25037), .C2(n5360), .ZN(n26131) );
  OAI22D0 U8944 ( .A1(n27143), .A2(n25038), .B1(n27142), .B2(n25039), .ZN(
        n26130) );
  OAI222D0 U8945 ( .A1(n24862), .A2(n25040), .B1(n25041), .B2(n5840), .C1(
        n25042), .C2(n5792), .ZN(n26129) );
  CKND0 U8946 ( .I(\Mem[44][26] ), .ZN(n24862) );
  AOI221D0 U8947 ( .A1(n27140), .A2(n25043), .B1(n27141), .B2(n25044), .C(
        n26133), .ZN(n26125) );
  OAI222D0 U8948 ( .A1(n25046), .A2(n6032), .B1(n24863), .B2(n25047), .C1(
        n25048), .C2(n4688), .ZN(n26133) );
  CKND0 U8949 ( .I(\Mem[45][26] ), .ZN(n24863) );
  NR4D0 U8950 ( .A1(n26134), .A2(n26135), .A3(n26136), .A4(n26137), .ZN(n26102) );
  OAI22D0 U8951 ( .A1(n25053), .A2(n5888), .B1(n25054), .B2(n5696), .ZN(n26137) );
  OAI222D0 U8952 ( .A1(n25055), .A2(n3824), .B1(n25056), .B2(n3872), .C1(
        n25057), .C2(n5936), .ZN(n26136) );
  OAI222D0 U8953 ( .A1(n25058), .A2(n3968), .B1(n25059), .B2(n4016), .C1(
        n25060), .C2(n3920), .ZN(n26135) );
  OAI222D0 U8954 ( .A1(n25061), .A2(n4112), .B1(n25062), .B2(n4160), .C1(
        n25063), .C2(n4064), .ZN(n26134) );
  NR4D0 U8955 ( .A1(n26138), .A2(n26139), .A3(n26140), .A4(n26141), .ZN(n26101) );
  OAI22D0 U8956 ( .A1(n25068), .A2(n2384), .B1(n25069), .B2(n2912), .ZN(n26141) );
  OAI222D0 U8957 ( .A1(n25070), .A2(n2480), .B1(n25071), .B2(n4304), .C1(
        n25072), .C2(n2624), .ZN(n26140) );
  OAI222D0 U8958 ( .A1(n25073), .A2(n4256), .B1(n24930), .B2(n3296), .C1(
        n25074), .C2(n4208), .ZN(n26139) );
  OAI222D0 U8959 ( .A1(n24932), .A2(n3392), .B1(n25075), .B2(n4832), .C1(
        n24931), .C2(n3344), .ZN(n26138) );
  ND4D0 U8960 ( .A1(n26142), .A2(n26143), .A3(n26144), .A4(n26145), .ZN(n2190)
         );
  AN4D0 U8961 ( .A1(n26146), .A2(n26147), .A3(n26148), .A4(n26149), .Z(n26145)
         );
  NR4D0 U8962 ( .A1(n26150), .A2(n26151), .A3(n26152), .A4(n26153), .ZN(n26149) );
  OAI222D0 U8963 ( .A1(n24979), .A2(n15557), .B1(n24980), .B2(n4447), .C1(
        n24964), .C2(n2239), .ZN(n26153) );
  OAI222D0 U8964 ( .A1(n24920), .A2(n2527), .B1(n24981), .B2(n5167), .C1(
        n24963), .C2(n2431), .ZN(n26152) );
  OAI222D0 U8965 ( .A1(n24982), .A2(n4927), .B1(n24983), .B2(n4975), .C1(
        n24984), .C2(n4879), .ZN(n26151) );
  OAI222D0 U8966 ( .A1(n24985), .A2(n4399), .B1(n24986), .B2(n3775), .C1(
        n24987), .C2(n4351), .ZN(n26150) );
  NR4D0 U8967 ( .A1(n26154), .A2(n26155), .A3(n26156), .A4(n26157), .ZN(n26148) );
  OAI22D0 U8968 ( .A1(n24922), .A2(n2815), .B1(n24992), .B2(n3727), .ZN(n26157) );
  OAI222D0 U8969 ( .A1(n24993), .A2(n18007), .B1(n24962), .B2(n2767), .C1(
        n24994), .C2(n18008), .ZN(n26156) );
  OAI222D0 U8970 ( .A1(n24995), .A2(n5215), .B1(n24961), .B2(n2671), .C1(
        n24921), .C2(n2719), .ZN(n26155) );
  OAI222D0 U8971 ( .A1(n24927), .A2(n3151), .B1(n24996), .B2(n4783), .C1(
        n24997), .C2(n15556), .ZN(n26154) );
  NR4D0 U8972 ( .A1(n26158), .A2(n26159), .A3(n26160), .A4(n26161), .ZN(n26147) );
  OAI22D0 U8973 ( .A1(n24928), .A2(n3199), .B1(n24926), .B2(n3103), .ZN(n26161) );
  OAI222D0 U8974 ( .A1(n25002), .A2(n3439), .B1(n24929), .B2(n3247), .C1(
        n24933), .C2(n2335), .ZN(n26160) );
  OAI222D0 U8975 ( .A1(n25003), .A2(n3583), .B1(n25004), .B2(n3487), .C1(
        n25005), .C2(n3535), .ZN(n26159) );
  OAI222D0 U8976 ( .A1(n24965), .A2(n2575), .B1(n25006), .B2(n3631), .C1(
        n25007), .C2(n3679), .ZN(n26158) );
  NR4D0 U8977 ( .A1(n26162), .A2(n26163), .A3(n26164), .A4(n26165), .ZN(n26146) );
  OAI22D0 U8978 ( .A1(n25012), .A2(n5119), .B1(n24966), .B2(n2287), .ZN(n26165) );
  OAI222D0 U8979 ( .A1(n24925), .A2(n3055), .B1(n24923), .B2(n2959), .C1(
        n24960), .C2(n2863), .ZN(n26164) );
  OAI222D0 U8980 ( .A1(n25013), .A2(n5503), .B1(n25014), .B2(n5551), .C1(
        n24924), .C2(n3007), .ZN(n26163) );
  OAI222D0 U8981 ( .A1(n25015), .A2(n6079), .B1(n25016), .B2(n5983), .C1(
        n25017), .C2(n6127), .ZN(n26162) );
  INR4D0 U8982 ( .A1(n26166), .B1(n26167), .B2(n26168), .B3(n26169), .ZN(
        n26144) );
  OAI222D0 U8983 ( .A1(n25022), .A2(n5455), .B1(n25023), .B2(n6319), .C1(
        n25024), .C2(n5407), .ZN(n26169) );
  OAI222D0 U8984 ( .A1(n25025), .A2(n4495), .B1(n25026), .B2(n24640), .C1(
        n25027), .C2(n5599), .ZN(n26168) );
  OR4D0 U8985 ( .A1(n26170), .A2(n26171), .A3(n26172), .A4(n26173), .Z(n26167)
         );
  OAI222D0 U8986 ( .A1(n25032), .A2(n4591), .B1(n25033), .B2(n5311), .C1(
        n25034), .C2(n6223), .ZN(n26173) );
  OAI222D0 U8987 ( .A1(n25035), .A2(n6175), .B1(n25036), .B2(n4543), .C1(
        n25037), .C2(n5359), .ZN(n26172) );
  OAI22D0 U8988 ( .A1(n27147), .A2(n25038), .B1(n27146), .B2(n25039), .ZN(
        n26171) );
  OAI222D0 U8989 ( .A1(n24860), .A2(n25040), .B1(n25041), .B2(n5839), .C1(
        n25042), .C2(n5791), .ZN(n26170) );
  CKND0 U8990 ( .I(\Mem[44][27] ), .ZN(n24860) );
  AOI221D0 U8991 ( .A1(n27144), .A2(n25043), .B1(n27145), .B2(n25044), .C(
        n26174), .ZN(n26166) );
  OAI222D0 U8992 ( .A1(n25046), .A2(n6031), .B1(n24861), .B2(n25047), .C1(
        n25048), .C2(n4687), .ZN(n26174) );
  CKND0 U8993 ( .I(\Mem[45][27] ), .ZN(n24861) );
  NR4D0 U8994 ( .A1(n26175), .A2(n26176), .A3(n26177), .A4(n26178), .ZN(n26143) );
  OAI22D0 U8995 ( .A1(n25053), .A2(n5887), .B1(n25054), .B2(n5695), .ZN(n26178) );
  OAI222D0 U8996 ( .A1(n25055), .A2(n3823), .B1(n25056), .B2(n3871), .C1(
        n25057), .C2(n5935), .ZN(n26177) );
  OAI222D0 U8997 ( .A1(n25058), .A2(n3967), .B1(n25059), .B2(n4015), .C1(
        n25060), .C2(n3919), .ZN(n26176) );
  OAI222D0 U8998 ( .A1(n25061), .A2(n4111), .B1(n25062), .B2(n4159), .C1(
        n25063), .C2(n4063), .ZN(n26175) );
  NR4D0 U8999 ( .A1(n26179), .A2(n26180), .A3(n26181), .A4(n26182), .ZN(n26142) );
  OAI22D0 U9000 ( .A1(n25068), .A2(n2383), .B1(n25069), .B2(n2911), .ZN(n26182) );
  OAI222D0 U9001 ( .A1(n25070), .A2(n2479), .B1(n25071), .B2(n4303), .C1(
        n25072), .C2(n2623), .ZN(n26181) );
  OAI222D0 U9002 ( .A1(n25073), .A2(n4255), .B1(n24930), .B2(n3295), .C1(
        n25074), .C2(n4207), .ZN(n26180) );
  OAI222D0 U9003 ( .A1(n24932), .A2(n3391), .B1(n25075), .B2(n4831), .C1(
        n24931), .C2(n3343), .ZN(n26179) );
  ND4D0 U9004 ( .A1(n26183), .A2(n26184), .A3(n26185), .A4(n26186), .ZN(n2189)
         );
  AN4D0 U9005 ( .A1(n26187), .A2(n26188), .A3(n26189), .A4(n26190), .Z(n26186)
         );
  NR4D0 U9006 ( .A1(n26191), .A2(n26192), .A3(n26193), .A4(n26194), .ZN(n26190) );
  OAI222D0 U9007 ( .A1(n24979), .A2(n15561), .B1(n24980), .B2(n4446), .C1(
        n24964), .C2(n2238), .ZN(n26194) );
  OAI222D0 U9008 ( .A1(n24920), .A2(n2526), .B1(n24981), .B2(n5166), .C1(
        n24963), .C2(n2430), .ZN(n26193) );
  OAI222D0 U9009 ( .A1(n24982), .A2(n4926), .B1(n24983), .B2(n4974), .C1(
        n24984), .C2(n4878), .ZN(n26192) );
  OAI222D0 U9010 ( .A1(n24985), .A2(n4398), .B1(n24986), .B2(n3774), .C1(
        n24987), .C2(n4350), .ZN(n26191) );
  NR4D0 U9011 ( .A1(n26195), .A2(n26196), .A3(n26197), .A4(n26198), .ZN(n26189) );
  OAI22D0 U9012 ( .A1(n24922), .A2(n2814), .B1(n24992), .B2(n3726), .ZN(n26198) );
  OAI222D0 U9013 ( .A1(n24993), .A2(n18010), .B1(n24962), .B2(n2766), .C1(
        n24994), .C2(n18011), .ZN(n26197) );
  OAI222D0 U9014 ( .A1(n24995), .A2(n5214), .B1(n24961), .B2(n2670), .C1(
        n24921), .C2(n2718), .ZN(n26196) );
  OAI222D0 U9015 ( .A1(n24927), .A2(n3150), .B1(n24996), .B2(n4782), .C1(
        n24997), .C2(n15560), .ZN(n26195) );
  NR4D0 U9016 ( .A1(n26199), .A2(n26200), .A3(n26201), .A4(n26202), .ZN(n26188) );
  OAI22D0 U9017 ( .A1(n24928), .A2(n3198), .B1(n24926), .B2(n3102), .ZN(n26202) );
  OAI222D0 U9018 ( .A1(n25002), .A2(n3438), .B1(n24929), .B2(n3246), .C1(
        n24933), .C2(n2334), .ZN(n26201) );
  OAI222D0 U9019 ( .A1(n25003), .A2(n3582), .B1(n25004), .B2(n3486), .C1(
        n25005), .C2(n3534), .ZN(n26200) );
  OAI222D0 U9020 ( .A1(n24965), .A2(n2574), .B1(n25006), .B2(n3630), .C1(
        n25007), .C2(n3678), .ZN(n26199) );
  NR4D0 U9021 ( .A1(n26203), .A2(n26204), .A3(n26205), .A4(n26206), .ZN(n26187) );
  OAI22D0 U9022 ( .A1(n25012), .A2(n5118), .B1(n24966), .B2(n2286), .ZN(n26206) );
  OAI222D0 U9023 ( .A1(n24925), .A2(n3054), .B1(n24923), .B2(n2958), .C1(
        n24960), .C2(n2862), .ZN(n26205) );
  OAI222D0 U9024 ( .A1(n25013), .A2(n5502), .B1(n25014), .B2(n5550), .C1(
        n24924), .C2(n3006), .ZN(n26204) );
  OAI222D0 U9025 ( .A1(n25015), .A2(n6078), .B1(n25016), .B2(n5982), .C1(
        n25017), .C2(n6126), .ZN(n26203) );
  INR4D0 U9026 ( .A1(n26207), .B1(n26208), .B2(n26209), .B3(n26210), .ZN(
        n26185) );
  OAI222D0 U9027 ( .A1(n25022), .A2(n5454), .B1(n25023), .B2(n6318), .C1(
        n25024), .C2(n5406), .ZN(n26210) );
  OAI222D0 U9028 ( .A1(n25025), .A2(n4494), .B1(n25026), .B2(n24643), .C1(
        n25027), .C2(n5598), .ZN(n26209) );
  OR4D0 U9029 ( .A1(n26211), .A2(n26212), .A3(n26213), .A4(n26214), .Z(n26208)
         );
  OAI222D0 U9030 ( .A1(n25032), .A2(n4590), .B1(n25033), .B2(n5310), .C1(
        n25034), .C2(n6222), .ZN(n26214) );
  OAI222D0 U9031 ( .A1(n25035), .A2(n6174), .B1(n25036), .B2(n4542), .C1(
        n25037), .C2(n5358), .ZN(n26213) );
  OAI22D0 U9032 ( .A1(n27151), .A2(n25038), .B1(n27150), .B2(n25039), .ZN(
        n26212) );
  OAI222D0 U9033 ( .A1(n24858), .A2(n25040), .B1(n25041), .B2(n5838), .C1(
        n25042), .C2(n5790), .ZN(n26211) );
  CKND0 U9034 ( .I(\Mem[44][28] ), .ZN(n24858) );
  AOI221D0 U9035 ( .A1(n27148), .A2(n25043), .B1(n27149), .B2(n25044), .C(
        n26215), .ZN(n26207) );
  OAI222D0 U9036 ( .A1(n25046), .A2(n6030), .B1(n24859), .B2(n25047), .C1(
        n25048), .C2(n4686), .ZN(n26215) );
  CKND0 U9037 ( .I(\Mem[45][28] ), .ZN(n24859) );
  NR4D0 U9038 ( .A1(n26216), .A2(n26217), .A3(n26218), .A4(n26219), .ZN(n26184) );
  OAI22D0 U9039 ( .A1(n25053), .A2(n5886), .B1(n25054), .B2(n5694), .ZN(n26219) );
  OAI222D0 U9040 ( .A1(n25055), .A2(n3822), .B1(n25056), .B2(n3870), .C1(
        n25057), .C2(n5934), .ZN(n26218) );
  OAI222D0 U9041 ( .A1(n25058), .A2(n3966), .B1(n25059), .B2(n4014), .C1(
        n25060), .C2(n3918), .ZN(n26217) );
  OAI222D0 U9042 ( .A1(n25061), .A2(n4110), .B1(n25062), .B2(n4158), .C1(
        n25063), .C2(n4062), .ZN(n26216) );
  NR4D0 U9043 ( .A1(n26220), .A2(n26221), .A3(n26222), .A4(n26223), .ZN(n26183) );
  OAI22D0 U9044 ( .A1(n25068), .A2(n2382), .B1(n25069), .B2(n2910), .ZN(n26223) );
  OAI222D0 U9045 ( .A1(n25070), .A2(n2478), .B1(n25071), .B2(n4302), .C1(
        n25072), .C2(n2622), .ZN(n26222) );
  OAI222D0 U9046 ( .A1(n25073), .A2(n4254), .B1(n24930), .B2(n3294), .C1(
        n25074), .C2(n4206), .ZN(n26221) );
  OAI222D0 U9047 ( .A1(n24932), .A2(n3390), .B1(n25075), .B2(n4830), .C1(
        n24931), .C2(n3342), .ZN(n26220) );
  ND4D0 U9048 ( .A1(n26224), .A2(n26225), .A3(n26226), .A4(n26227), .ZN(n2188)
         );
  AN4D0 U9049 ( .A1(n26228), .A2(n26229), .A3(n26230), .A4(n26231), .Z(n26227)
         );
  NR4D0 U9050 ( .A1(n26232), .A2(n26233), .A3(n26234), .A4(n26235), .ZN(n26231) );
  OAI222D0 U9051 ( .A1(n24979), .A2(n15565), .B1(n24980), .B2(n4445), .C1(
        n24964), .C2(n2237), .ZN(n26235) );
  OAI222D0 U9052 ( .A1(n24920), .A2(n2525), .B1(n24981), .B2(n5165), .C1(
        n24963), .C2(n2429), .ZN(n26234) );
  OAI222D0 U9053 ( .A1(n24982), .A2(n4925), .B1(n24983), .B2(n4973), .C1(
        n24984), .C2(n4877), .ZN(n26233) );
  OAI222D0 U9054 ( .A1(n24985), .A2(n4397), .B1(n24986), .B2(n3773), .C1(
        n24987), .C2(n4349), .ZN(n26232) );
  NR4D0 U9055 ( .A1(n26236), .A2(n26237), .A3(n26238), .A4(n26239), .ZN(n26230) );
  OAI22D0 U9056 ( .A1(n24922), .A2(n2813), .B1(n24992), .B2(n3725), .ZN(n26239) );
  OAI222D0 U9057 ( .A1(n24993), .A2(n18013), .B1(n24962), .B2(n2765), .C1(
        n24994), .C2(n18014), .ZN(n26238) );
  OAI222D0 U9058 ( .A1(n24995), .A2(n5213), .B1(n24961), .B2(n2669), .C1(
        n24921), .C2(n2717), .ZN(n26237) );
  OAI222D0 U9059 ( .A1(n24927), .A2(n3149), .B1(n24996), .B2(n4781), .C1(
        n24997), .C2(n15564), .ZN(n26236) );
  NR4D0 U9060 ( .A1(n26240), .A2(n26241), .A3(n26242), .A4(n26243), .ZN(n26229) );
  OAI22D0 U9061 ( .A1(n24928), .A2(n3197), .B1(n24926), .B2(n3101), .ZN(n26243) );
  OAI222D0 U9062 ( .A1(n25002), .A2(n3437), .B1(n24929), .B2(n3245), .C1(
        n24933), .C2(n2333), .ZN(n26242) );
  OAI222D0 U9063 ( .A1(n25003), .A2(n3581), .B1(n25004), .B2(n3485), .C1(
        n25005), .C2(n3533), .ZN(n26241) );
  OAI222D0 U9064 ( .A1(n24965), .A2(n2573), .B1(n25006), .B2(n3629), .C1(
        n25007), .C2(n3677), .ZN(n26240) );
  NR4D0 U9065 ( .A1(n26244), .A2(n26245), .A3(n26246), .A4(n26247), .ZN(n26228) );
  OAI22D0 U9066 ( .A1(n25012), .A2(n5117), .B1(n24966), .B2(n2285), .ZN(n26247) );
  OAI222D0 U9067 ( .A1(n24925), .A2(n3053), .B1(n24923), .B2(n2957), .C1(
        n24960), .C2(n2861), .ZN(n26246) );
  OAI222D0 U9068 ( .A1(n25013), .A2(n5501), .B1(n25014), .B2(n5549), .C1(
        n24924), .C2(n3005), .ZN(n26245) );
  OAI222D0 U9069 ( .A1(n25015), .A2(n6077), .B1(n25016), .B2(n5981), .C1(
        n25017), .C2(n6125), .ZN(n26244) );
  INR4D0 U9070 ( .A1(n26248), .B1(n26249), .B2(n26250), .B3(n26251), .ZN(
        n26226) );
  OAI222D0 U9071 ( .A1(n25022), .A2(n5453), .B1(n25023), .B2(n6317), .C1(
        n25024), .C2(n5405), .ZN(n26251) );
  OAI222D0 U9072 ( .A1(n25025), .A2(n4493), .B1(n25026), .B2(n24646), .C1(
        n25027), .C2(n5597), .ZN(n26250) );
  OR4D0 U9073 ( .A1(n26252), .A2(n26253), .A3(n26254), .A4(n26255), .Z(n26249)
         );
  OAI222D0 U9074 ( .A1(n25032), .A2(n4589), .B1(n25033), .B2(n5309), .C1(
        n25034), .C2(n6221), .ZN(n26255) );
  OAI222D0 U9075 ( .A1(n25035), .A2(n6173), .B1(n25036), .B2(n4541), .C1(
        n25037), .C2(n5357), .ZN(n26254) );
  OAI22D0 U9076 ( .A1(n27155), .A2(n25038), .B1(n27154), .B2(n25039), .ZN(
        n26253) );
  OAI222D0 U9077 ( .A1(n24856), .A2(n25040), .B1(n25041), .B2(n5837), .C1(
        n25042), .C2(n5789), .ZN(n26252) );
  CKND0 U9078 ( .I(\Mem[44][29] ), .ZN(n24856) );
  AOI221D0 U9079 ( .A1(n27152), .A2(n25043), .B1(n27153), .B2(n25044), .C(
        n26256), .ZN(n26248) );
  OAI222D0 U9080 ( .A1(n25046), .A2(n6029), .B1(n24857), .B2(n25047), .C1(
        n25048), .C2(n4685), .ZN(n26256) );
  CKND0 U9081 ( .I(\Mem[45][29] ), .ZN(n24857) );
  NR4D0 U9082 ( .A1(n26257), .A2(n26258), .A3(n26259), .A4(n26260), .ZN(n26225) );
  OAI22D0 U9083 ( .A1(n25053), .A2(n5885), .B1(n25054), .B2(n5693), .ZN(n26260) );
  OAI222D0 U9084 ( .A1(n25055), .A2(n3821), .B1(n25056), .B2(n3869), .C1(
        n25057), .C2(n5933), .ZN(n26259) );
  OAI222D0 U9085 ( .A1(n25058), .A2(n3965), .B1(n25059), .B2(n4013), .C1(
        n25060), .C2(n3917), .ZN(n26258) );
  OAI222D0 U9086 ( .A1(n25061), .A2(n4109), .B1(n25062), .B2(n4157), .C1(
        n25063), .C2(n4061), .ZN(n26257) );
  NR4D0 U9087 ( .A1(n26261), .A2(n26262), .A3(n26263), .A4(n26264), .ZN(n26224) );
  OAI22D0 U9088 ( .A1(n25068), .A2(n2381), .B1(n25069), .B2(n2909), .ZN(n26264) );
  OAI222D0 U9089 ( .A1(n25070), .A2(n2477), .B1(n25071), .B2(n4301), .C1(
        n25072), .C2(n2621), .ZN(n26263) );
  OAI222D0 U9090 ( .A1(n25073), .A2(n4253), .B1(n24930), .B2(n3293), .C1(
        n25074), .C2(n4205), .ZN(n26262) );
  OAI222D0 U9091 ( .A1(n24932), .A2(n3389), .B1(n25075), .B2(n4829), .C1(
        n24931), .C2(n3341), .ZN(n26261) );
  ND4D0 U9092 ( .A1(n26265), .A2(n26266), .A3(n26267), .A4(n26268), .ZN(n2187)
         );
  AN4D0 U9093 ( .A1(n26269), .A2(n26270), .A3(n26271), .A4(n26272), .Z(n26268)
         );
  NR4D0 U9094 ( .A1(n26273), .A2(n26274), .A3(n26275), .A4(n26276), .ZN(n26272) );
  OAI222D0 U9095 ( .A1(n24979), .A2(n15569), .B1(n24980), .B2(n4444), .C1(
        n24964), .C2(n2236), .ZN(n26276) );
  OAI222D0 U9096 ( .A1(n24920), .A2(n2524), .B1(n24981), .B2(n5164), .C1(
        n24963), .C2(n2428), .ZN(n26275) );
  OAI222D0 U9097 ( .A1(n24982), .A2(n4924), .B1(n24983), .B2(n4972), .C1(
        n24984), .C2(n4876), .ZN(n26274) );
  OAI222D0 U9098 ( .A1(n24985), .A2(n4396), .B1(n24986), .B2(n3772), .C1(
        n24987), .C2(n4348), .ZN(n26273) );
  NR4D0 U9099 ( .A1(n26277), .A2(n26278), .A3(n26279), .A4(n26280), .ZN(n26271) );
  OAI22D0 U9100 ( .A1(n24922), .A2(n2812), .B1(n24992), .B2(n3724), .ZN(n26280) );
  OAI222D0 U9101 ( .A1(n24993), .A2(n18016), .B1(n24962), .B2(n2764), .C1(
        n24994), .C2(n18017), .ZN(n26279) );
  OAI222D0 U9102 ( .A1(n24995), .A2(n5212), .B1(n24961), .B2(n2668), .C1(
        n24921), .C2(n2716), .ZN(n26278) );
  OAI222D0 U9103 ( .A1(n24927), .A2(n3148), .B1(n24996), .B2(n4780), .C1(
        n24997), .C2(n15568), .ZN(n26277) );
  NR4D0 U9104 ( .A1(n26281), .A2(n26282), .A3(n26283), .A4(n26284), .ZN(n26270) );
  OAI22D0 U9105 ( .A1(n24928), .A2(n3196), .B1(n24926), .B2(n3100), .ZN(n26284) );
  OAI222D0 U9106 ( .A1(n25002), .A2(n3436), .B1(n24929), .B2(n3244), .C1(
        n24933), .C2(n2332), .ZN(n26283) );
  OAI222D0 U9107 ( .A1(n25003), .A2(n3580), .B1(n25004), .B2(n3484), .C1(
        n25005), .C2(n3532), .ZN(n26282) );
  OAI222D0 U9108 ( .A1(n24965), .A2(n2572), .B1(n25006), .B2(n3628), .C1(
        n25007), .C2(n3676), .ZN(n26281) );
  NR4D0 U9109 ( .A1(n26285), .A2(n26286), .A3(n26287), .A4(n26288), .ZN(n26269) );
  OAI22D0 U9110 ( .A1(n25012), .A2(n5116), .B1(n24966), .B2(n2284), .ZN(n26288) );
  OAI222D0 U9111 ( .A1(n24925), .A2(n3052), .B1(n24923), .B2(n2956), .C1(
        n24960), .C2(n2860), .ZN(n26287) );
  OAI222D0 U9112 ( .A1(n25013), .A2(n5500), .B1(n25014), .B2(n5548), .C1(
        n24924), .C2(n3004), .ZN(n26286) );
  OAI222D0 U9113 ( .A1(n25015), .A2(n6076), .B1(n25016), .B2(n5980), .C1(
        n25017), .C2(n6124), .ZN(n26285) );
  INR4D0 U9114 ( .A1(n26289), .B1(n26290), .B2(n26291), .B3(n26292), .ZN(
        n26267) );
  OAI222D0 U9115 ( .A1(n25022), .A2(n5452), .B1(n25023), .B2(n6316), .C1(
        n25024), .C2(n5404), .ZN(n26292) );
  OAI222D0 U9116 ( .A1(n25025), .A2(n4492), .B1(n25026), .B2(n24649), .C1(
        n25027), .C2(n5596), .ZN(n26291) );
  OR4D0 U9117 ( .A1(n26293), .A2(n26294), .A3(n26295), .A4(n26296), .Z(n26290)
         );
  OAI222D0 U9118 ( .A1(n25032), .A2(n4588), .B1(n25033), .B2(n5308), .C1(
        n25034), .C2(n6220), .ZN(n26296) );
  OAI222D0 U9119 ( .A1(n25035), .A2(n6172), .B1(n25036), .B2(n4540), .C1(
        n25037), .C2(n5356), .ZN(n26295) );
  OAI22D0 U9120 ( .A1(n27159), .A2(n25038), .B1(n27158), .B2(n25039), .ZN(
        n26294) );
  OAI222D0 U9121 ( .A1(n24854), .A2(n25040), .B1(n25041), .B2(n5836), .C1(
        n25042), .C2(n5788), .ZN(n26293) );
  CKND0 U9122 ( .I(\Mem[44][30] ), .ZN(n24854) );
  AOI221D0 U9123 ( .A1(n27156), .A2(n25043), .B1(n27157), .B2(n25044), .C(
        n26297), .ZN(n26289) );
  OAI222D0 U9124 ( .A1(n25046), .A2(n6028), .B1(n24855), .B2(n25047), .C1(
        n25048), .C2(n4684), .ZN(n26297) );
  CKND0 U9125 ( .I(\Mem[45][30] ), .ZN(n24855) );
  NR4D0 U9126 ( .A1(n26298), .A2(n26299), .A3(n26300), .A4(n26301), .ZN(n26266) );
  OAI22D0 U9127 ( .A1(n25053), .A2(n5884), .B1(n25054), .B2(n5692), .ZN(n26301) );
  OAI222D0 U9128 ( .A1(n25055), .A2(n3820), .B1(n25056), .B2(n3868), .C1(
        n25057), .C2(n5932), .ZN(n26300) );
  OAI222D0 U9129 ( .A1(n25058), .A2(n3964), .B1(n25059), .B2(n4012), .C1(
        n25060), .C2(n3916), .ZN(n26299) );
  OAI222D0 U9130 ( .A1(n25061), .A2(n4108), .B1(n25062), .B2(n4156), .C1(
        n25063), .C2(n4060), .ZN(n26298) );
  NR4D0 U9131 ( .A1(n26302), .A2(n26303), .A3(n26304), .A4(n26305), .ZN(n26265) );
  OAI22D0 U9132 ( .A1(n25068), .A2(n2380), .B1(n25069), .B2(n2908), .ZN(n26305) );
  OAI222D0 U9133 ( .A1(n25070), .A2(n2476), .B1(n25071), .B2(n4300), .C1(
        n25072), .C2(n2620), .ZN(n26304) );
  OAI222D0 U9134 ( .A1(n25073), .A2(n4252), .B1(n24930), .B2(n3292), .C1(
        n25074), .C2(n4204), .ZN(n26303) );
  OAI222D0 U9135 ( .A1(n24932), .A2(n3388), .B1(n25075), .B2(n4828), .C1(
        n24931), .C2(n3340), .ZN(n26302) );
  ND4D0 U9136 ( .A1(n26306), .A2(n26307), .A3(n26308), .A4(n26309), .ZN(n2186)
         );
  AN4D0 U9137 ( .A1(n26310), .A2(n26311), .A3(n26312), .A4(n26313), .Z(n26309)
         );
  NR4D0 U9138 ( .A1(n26314), .A2(n26315), .A3(n26316), .A4(n26317), .ZN(n26313) );
  OAI222D0 U9139 ( .A1(n24979), .A2(n15573), .B1(n24980), .B2(n4443), .C1(
        n24964), .C2(n2235), .ZN(n26317) );
  OAI222D0 U9140 ( .A1(n24920), .A2(n2523), .B1(n24981), .B2(n5163), .C1(
        n24963), .C2(n2427), .ZN(n26316) );
  OAI222D0 U9141 ( .A1(n24982), .A2(n4923), .B1(n24983), .B2(n4971), .C1(
        n24984), .C2(n4875), .ZN(n26315) );
  OAI222D0 U9142 ( .A1(n24985), .A2(n4395), .B1(n24986), .B2(n3771), .C1(
        n24987), .C2(n4347), .ZN(n26314) );
  NR4D0 U9143 ( .A1(n26318), .A2(n26319), .A3(n26320), .A4(n26321), .ZN(n26312) );
  OAI22D0 U9144 ( .A1(n24922), .A2(n2811), .B1(n24992), .B2(n3723), .ZN(n26321) );
  OAI222D0 U9145 ( .A1(n24993), .A2(n18019), .B1(n24962), .B2(n2763), .C1(
        n24994), .C2(n18020), .ZN(n26320) );
  OAI222D0 U9146 ( .A1(n24995), .A2(n5211), .B1(n24961), .B2(n2667), .C1(
        n24921), .C2(n2715), .ZN(n26319) );
  OAI222D0 U9147 ( .A1(n24927), .A2(n3147), .B1(n24996), .B2(n4779), .C1(
        n24997), .C2(n15572), .ZN(n26318) );
  NR4D0 U9148 ( .A1(n26322), .A2(n26323), .A3(n26324), .A4(n26325), .ZN(n26311) );
  OAI22D0 U9149 ( .A1(n24928), .A2(n3195), .B1(n24926), .B2(n3099), .ZN(n26325) );
  OAI222D0 U9150 ( .A1(n25002), .A2(n3435), .B1(n24929), .B2(n3243), .C1(
        n24933), .C2(n2331), .ZN(n26324) );
  OAI222D0 U9151 ( .A1(n25003), .A2(n3579), .B1(n25004), .B2(n3483), .C1(
        n25005), .C2(n3531), .ZN(n26323) );
  OAI222D0 U9152 ( .A1(n24965), .A2(n2571), .B1(n25006), .B2(n3627), .C1(
        n25007), .C2(n3675), .ZN(n26322) );
  NR4D0 U9153 ( .A1(n26326), .A2(n26327), .A3(n26328), .A4(n26329), .ZN(n26310) );
  OAI22D0 U9154 ( .A1(n25012), .A2(n5115), .B1(n24966), .B2(n2283), .ZN(n26329) );
  OAI222D0 U9155 ( .A1(n24925), .A2(n3051), .B1(n24923), .B2(n2955), .C1(
        n24960), .C2(n2859), .ZN(n26328) );
  OAI222D0 U9156 ( .A1(n25013), .A2(n5499), .B1(n25014), .B2(n5547), .C1(
        n24924), .C2(n3003), .ZN(n26327) );
  OAI222D0 U9157 ( .A1(n25015), .A2(n6075), .B1(n25016), .B2(n5979), .C1(
        n25017), .C2(n6123), .ZN(n26326) );
  INR4D0 U9158 ( .A1(n26330), .B1(n26331), .B2(n26332), .B3(n26333), .ZN(
        n26308) );
  OAI222D0 U9159 ( .A1(n25022), .A2(n5451), .B1(n25023), .B2(n6315), .C1(
        n25024), .C2(n5403), .ZN(n26333) );
  OAI222D0 U9160 ( .A1(n25025), .A2(n4491), .B1(n25026), .B2(n24652), .C1(
        n25027), .C2(n5595), .ZN(n26332) );
  OR4D0 U9161 ( .A1(n26334), .A2(n26335), .A3(n26336), .A4(n26337), .Z(n26331)
         );
  OAI222D0 U9162 ( .A1(n25032), .A2(n4587), .B1(n25033), .B2(n5307), .C1(
        n25034), .C2(n6219), .ZN(n26337) );
  OAI222D0 U9163 ( .A1(n25035), .A2(n6171), .B1(n25036), .B2(n4539), .C1(
        n25037), .C2(n5355), .ZN(n26336) );
  OAI22D0 U9164 ( .A1(n27163), .A2(n25038), .B1(n27162), .B2(n25039), .ZN(
        n26335) );
  OAI222D0 U9165 ( .A1(n24852), .A2(n25040), .B1(n25041), .B2(n5835), .C1(
        n25042), .C2(n5787), .ZN(n26334) );
  CKND0 U9166 ( .I(\Mem[44][31] ), .ZN(n24852) );
  AOI221D0 U9167 ( .A1(n27160), .A2(n25043), .B1(n27161), .B2(n25044), .C(
        n26338), .ZN(n26330) );
  OAI222D0 U9168 ( .A1(n25046), .A2(n6027), .B1(n24853), .B2(n25047), .C1(
        n25048), .C2(n4683), .ZN(n26338) );
  CKND0 U9169 ( .I(\Mem[45][31] ), .ZN(n24853) );
  NR4D0 U9170 ( .A1(n26339), .A2(n26340), .A3(n26341), .A4(n26342), .ZN(n26307) );
  OAI22D0 U9171 ( .A1(n25053), .A2(n5883), .B1(n25054), .B2(n5691), .ZN(n26342) );
  OAI222D0 U9172 ( .A1(n25055), .A2(n3819), .B1(n25056), .B2(n3867), .C1(
        n25057), .C2(n5931), .ZN(n26341) );
  OAI222D0 U9173 ( .A1(n25058), .A2(n3963), .B1(n25059), .B2(n4011), .C1(
        n25060), .C2(n3915), .ZN(n26340) );
  OAI222D0 U9174 ( .A1(n25061), .A2(n4107), .B1(n25062), .B2(n4155), .C1(
        n25063), .C2(n4059), .ZN(n26339) );
  NR4D0 U9175 ( .A1(n26343), .A2(n26344), .A3(n26345), .A4(n26346), .ZN(n26306) );
  OAI22D0 U9176 ( .A1(n25068), .A2(n2379), .B1(n25069), .B2(n2907), .ZN(n26346) );
  OAI222D0 U9177 ( .A1(n25070), .A2(n2475), .B1(n25071), .B2(n4299), .C1(
        n25072), .C2(n2619), .ZN(n26345) );
  OAI222D0 U9178 ( .A1(n25073), .A2(n4251), .B1(n24930), .B2(n3291), .C1(
        n25074), .C2(n4203), .ZN(n26344) );
  OAI222D0 U9179 ( .A1(n24932), .A2(n3387), .B1(n25075), .B2(n4827), .C1(
        n24931), .C2(n3339), .ZN(n26343) );
  ND4D0 U9180 ( .A1(n26347), .A2(n26348), .A3(n26349), .A4(n26350), .ZN(n2185)
         );
  AN4D0 U9181 ( .A1(n26351), .A2(n26352), .A3(n26353), .A4(n26354), .Z(n26350)
         );
  NR4D0 U9182 ( .A1(n26355), .A2(n26356), .A3(n26357), .A4(n26358), .ZN(n26354) );
  OAI222D0 U9183 ( .A1(n24979), .A2(n15577), .B1(n24980), .B2(n4442), .C1(
        n24964), .C2(n2234), .ZN(n26358) );
  OAI222D0 U9184 ( .A1(n24920), .A2(n2522), .B1(n24981), .B2(n5162), .C1(
        n24963), .C2(n2426), .ZN(n26357) );
  OAI222D0 U9185 ( .A1(n24982), .A2(n4922), .B1(n24983), .B2(n4970), .C1(
        n24984), .C2(n4874), .ZN(n26356) );
  OAI222D0 U9186 ( .A1(n24985), .A2(n4394), .B1(n24986), .B2(n3770), .C1(
        n24987), .C2(n4346), .ZN(n26355) );
  NR4D0 U9187 ( .A1(n26359), .A2(n26360), .A3(n26361), .A4(n26362), .ZN(n26353) );
  OAI22D0 U9188 ( .A1(n24922), .A2(n2810), .B1(n24992), .B2(n3722), .ZN(n26362) );
  OAI222D0 U9189 ( .A1(n24993), .A2(n18022), .B1(n24962), .B2(n2762), .C1(
        n24994), .C2(n18023), .ZN(n26361) );
  OAI222D0 U9190 ( .A1(n24995), .A2(n5210), .B1(n24961), .B2(n2666), .C1(
        n24921), .C2(n2714), .ZN(n26360) );
  OAI222D0 U9191 ( .A1(n24927), .A2(n3146), .B1(n24996), .B2(n4778), .C1(
        n24997), .C2(n15576), .ZN(n26359) );
  NR4D0 U9192 ( .A1(n26363), .A2(n26364), .A3(n26365), .A4(n26366), .ZN(n26352) );
  OAI22D0 U9193 ( .A1(n24928), .A2(n3194), .B1(n24926), .B2(n3098), .ZN(n26366) );
  OAI222D0 U9194 ( .A1(n25002), .A2(n3434), .B1(n24929), .B2(n3242), .C1(
        n24933), .C2(n2330), .ZN(n26365) );
  OAI222D0 U9195 ( .A1(n25003), .A2(n3578), .B1(n25004), .B2(n3482), .C1(
        n25005), .C2(n3530), .ZN(n26364) );
  OAI222D0 U9196 ( .A1(n24965), .A2(n2570), .B1(n25006), .B2(n3626), .C1(
        n25007), .C2(n3674), .ZN(n26363) );
  NR4D0 U9197 ( .A1(n26367), .A2(n26368), .A3(n26369), .A4(n26370), .ZN(n26351) );
  OAI22D0 U9198 ( .A1(n25012), .A2(n5114), .B1(n24966), .B2(n2282), .ZN(n26370) );
  OAI222D0 U9199 ( .A1(n24925), .A2(n3050), .B1(n24923), .B2(n2954), .C1(
        n24960), .C2(n2858), .ZN(n26369) );
  OAI222D0 U9200 ( .A1(n25013), .A2(n5498), .B1(n25014), .B2(n5546), .C1(
        n24924), .C2(n3002), .ZN(n26368) );
  OAI222D0 U9201 ( .A1(n25015), .A2(n6074), .B1(n25016), .B2(n5978), .C1(
        n25017), .C2(n6122), .ZN(n26367) );
  INR4D0 U9202 ( .A1(n26371), .B1(n26372), .B2(n26373), .B3(n26374), .ZN(
        n26349) );
  OAI222D0 U9203 ( .A1(n25022), .A2(n5450), .B1(n25023), .B2(n6314), .C1(
        n25024), .C2(n5402), .ZN(n26374) );
  OAI222D0 U9204 ( .A1(n25025), .A2(n4490), .B1(n25026), .B2(n24655), .C1(
        n25027), .C2(n5594), .ZN(n26373) );
  OR4D0 U9205 ( .A1(n26375), .A2(n26376), .A3(n26377), .A4(n26378), .Z(n26372)
         );
  OAI222D0 U9206 ( .A1(n25032), .A2(n4586), .B1(n25033), .B2(n5306), .C1(
        n25034), .C2(n6218), .ZN(n26378) );
  OAI222D0 U9207 ( .A1(n25035), .A2(n6170), .B1(n25036), .B2(n4538), .C1(
        n25037), .C2(n5354), .ZN(n26377) );
  OAI22D0 U9208 ( .A1(n27167), .A2(n25038), .B1(n27166), .B2(n25039), .ZN(
        n26376) );
  OAI222D0 U9209 ( .A1(n24850), .A2(n25040), .B1(n25041), .B2(n5834), .C1(
        n25042), .C2(n5786), .ZN(n26375) );
  CKND0 U9210 ( .I(\Mem[44][32] ), .ZN(n24850) );
  AOI221D0 U9211 ( .A1(n27164), .A2(n25043), .B1(n27165), .B2(n25044), .C(
        n26379), .ZN(n26371) );
  OAI222D0 U9212 ( .A1(n25046), .A2(n6026), .B1(n24851), .B2(n25047), .C1(
        n25048), .C2(n4682), .ZN(n26379) );
  CKND0 U9213 ( .I(\Mem[45][32] ), .ZN(n24851) );
  NR4D0 U9214 ( .A1(n26380), .A2(n26381), .A3(n26382), .A4(n26383), .ZN(n26348) );
  OAI22D0 U9215 ( .A1(n25053), .A2(n5882), .B1(n25054), .B2(n5690), .ZN(n26383) );
  OAI222D0 U9216 ( .A1(n25055), .A2(n3818), .B1(n25056), .B2(n3866), .C1(
        n25057), .C2(n5930), .ZN(n26382) );
  OAI222D0 U9217 ( .A1(n25058), .A2(n3962), .B1(n25059), .B2(n4010), .C1(
        n25060), .C2(n3914), .ZN(n26381) );
  OAI222D0 U9218 ( .A1(n25061), .A2(n4106), .B1(n25062), .B2(n4154), .C1(
        n25063), .C2(n4058), .ZN(n26380) );
  NR4D0 U9219 ( .A1(n26384), .A2(n26385), .A3(n26386), .A4(n26387), .ZN(n26347) );
  OAI22D0 U9220 ( .A1(n25068), .A2(n2378), .B1(n25069), .B2(n2906), .ZN(n26387) );
  OAI222D0 U9221 ( .A1(n25070), .A2(n2474), .B1(n25071), .B2(n4298), .C1(
        n25072), .C2(n2618), .ZN(n26386) );
  OAI222D0 U9222 ( .A1(n25073), .A2(n4250), .B1(n24930), .B2(n3290), .C1(
        n25074), .C2(n4202), .ZN(n26385) );
  OAI222D0 U9223 ( .A1(n24932), .A2(n3386), .B1(n25075), .B2(n4826), .C1(
        n24931), .C2(n3338), .ZN(n26384) );
  ND4D0 U9224 ( .A1(n26388), .A2(n26389), .A3(n26390), .A4(n26391), .ZN(n2184)
         );
  AN4D0 U9225 ( .A1(n26392), .A2(n26393), .A3(n26394), .A4(n26395), .Z(n26391)
         );
  NR4D0 U9226 ( .A1(n26396), .A2(n26397), .A3(n26398), .A4(n26399), .ZN(n26395) );
  OAI222D0 U9227 ( .A1(n24979), .A2(n15581), .B1(n24980), .B2(n4441), .C1(
        n24964), .C2(n2233), .ZN(n26399) );
  OAI222D0 U9228 ( .A1(n24920), .A2(n2521), .B1(n24981), .B2(n5161), .C1(
        n24963), .C2(n2425), .ZN(n26398) );
  OAI222D0 U9229 ( .A1(n24982), .A2(n4921), .B1(n24983), .B2(n4969), .C1(
        n24984), .C2(n4873), .ZN(n26397) );
  OAI222D0 U9230 ( .A1(n24985), .A2(n4393), .B1(n24986), .B2(n3769), .C1(
        n24987), .C2(n4345), .ZN(n26396) );
  NR4D0 U9231 ( .A1(n26400), .A2(n26401), .A3(n26402), .A4(n26403), .ZN(n26394) );
  OAI22D0 U9232 ( .A1(n24922), .A2(n2809), .B1(n24992), .B2(n3721), .ZN(n26403) );
  OAI222D0 U9233 ( .A1(n24993), .A2(n18025), .B1(n24962), .B2(n2761), .C1(
        n24994), .C2(n18026), .ZN(n26402) );
  OAI222D0 U9234 ( .A1(n24995), .A2(n5209), .B1(n24961), .B2(n2665), .C1(
        n24921), .C2(n2713), .ZN(n26401) );
  OAI222D0 U9235 ( .A1(n24927), .A2(n3145), .B1(n24996), .B2(n4777), .C1(
        n24997), .C2(n15580), .ZN(n26400) );
  NR4D0 U9236 ( .A1(n26404), .A2(n26405), .A3(n26406), .A4(n26407), .ZN(n26393) );
  OAI22D0 U9237 ( .A1(n24928), .A2(n3193), .B1(n24926), .B2(n3097), .ZN(n26407) );
  OAI222D0 U9238 ( .A1(n25002), .A2(n3433), .B1(n24929), .B2(n3241), .C1(
        n24933), .C2(n2329), .ZN(n26406) );
  OAI222D0 U9239 ( .A1(n25003), .A2(n3577), .B1(n25004), .B2(n3481), .C1(
        n25005), .C2(n3529), .ZN(n26405) );
  OAI222D0 U9240 ( .A1(n24965), .A2(n2569), .B1(n25006), .B2(n3625), .C1(
        n25007), .C2(n3673), .ZN(n26404) );
  NR4D0 U9241 ( .A1(n26408), .A2(n26409), .A3(n26410), .A4(n26411), .ZN(n26392) );
  OAI22D0 U9242 ( .A1(n25012), .A2(n5113), .B1(n24966), .B2(n2281), .ZN(n26411) );
  OAI222D0 U9243 ( .A1(n24925), .A2(n3049), .B1(n24923), .B2(n2953), .C1(
        n24960), .C2(n2857), .ZN(n26410) );
  OAI222D0 U9244 ( .A1(n25013), .A2(n5497), .B1(n25014), .B2(n5545), .C1(
        n24924), .C2(n3001), .ZN(n26409) );
  OAI222D0 U9245 ( .A1(n25015), .A2(n6073), .B1(n25016), .B2(n5977), .C1(
        n25017), .C2(n6121), .ZN(n26408) );
  INR4D0 U9246 ( .A1(n26412), .B1(n26413), .B2(n26414), .B3(n26415), .ZN(
        n26390) );
  OAI222D0 U9247 ( .A1(n25022), .A2(n5449), .B1(n25023), .B2(n6313), .C1(
        n25024), .C2(n5401), .ZN(n26415) );
  OAI222D0 U9248 ( .A1(n25025), .A2(n4489), .B1(n25026), .B2(n24658), .C1(
        n25027), .C2(n5593), .ZN(n26414) );
  OR4D0 U9249 ( .A1(n26416), .A2(n26417), .A3(n26418), .A4(n26419), .Z(n26413)
         );
  OAI222D0 U9250 ( .A1(n25032), .A2(n4585), .B1(n25033), .B2(n5305), .C1(
        n25034), .C2(n6217), .ZN(n26419) );
  OAI222D0 U9251 ( .A1(n25035), .A2(n6169), .B1(n25036), .B2(n4537), .C1(
        n25037), .C2(n5353), .ZN(n26418) );
  OAI22D0 U9252 ( .A1(n27171), .A2(n25038), .B1(n27170), .B2(n25039), .ZN(
        n26417) );
  OAI222D0 U9253 ( .A1(n24848), .A2(n25040), .B1(n25041), .B2(n5833), .C1(
        n25042), .C2(n5785), .ZN(n26416) );
  CKND0 U9254 ( .I(\Mem[44][33] ), .ZN(n24848) );
  AOI221D0 U9255 ( .A1(n27168), .A2(n25043), .B1(n27169), .B2(n25044), .C(
        n26420), .ZN(n26412) );
  OAI222D0 U9256 ( .A1(n25046), .A2(n6025), .B1(n24849), .B2(n25047), .C1(
        n25048), .C2(n4681), .ZN(n26420) );
  CKND0 U9257 ( .I(\Mem[45][33] ), .ZN(n24849) );
  NR4D0 U9258 ( .A1(n26421), .A2(n26422), .A3(n26423), .A4(n26424), .ZN(n26389) );
  OAI22D0 U9259 ( .A1(n25053), .A2(n5881), .B1(n25054), .B2(n5689), .ZN(n26424) );
  OAI222D0 U9260 ( .A1(n25055), .A2(n3817), .B1(n25056), .B2(n3865), .C1(
        n25057), .C2(n5929), .ZN(n26423) );
  OAI222D0 U9261 ( .A1(n25058), .A2(n3961), .B1(n25059), .B2(n4009), .C1(
        n25060), .C2(n3913), .ZN(n26422) );
  OAI222D0 U9262 ( .A1(n25061), .A2(n4105), .B1(n25062), .B2(n4153), .C1(
        n25063), .C2(n4057), .ZN(n26421) );
  NR4D0 U9263 ( .A1(n26425), .A2(n26426), .A3(n26427), .A4(n26428), .ZN(n26388) );
  OAI22D0 U9264 ( .A1(n25068), .A2(n2377), .B1(n25069), .B2(n2905), .ZN(n26428) );
  OAI222D0 U9265 ( .A1(n25070), .A2(n2473), .B1(n25071), .B2(n4297), .C1(
        n25072), .C2(n2617), .ZN(n26427) );
  OAI222D0 U9266 ( .A1(n25073), .A2(n4249), .B1(n24930), .B2(n3289), .C1(
        n25074), .C2(n4201), .ZN(n26426) );
  OAI222D0 U9267 ( .A1(n24932), .A2(n3385), .B1(n25075), .B2(n4825), .C1(
        n24931), .C2(n3337), .ZN(n26425) );
  ND4D0 U9268 ( .A1(n26429), .A2(n26430), .A3(n26431), .A4(n26432), .ZN(n2183)
         );
  AN4D0 U9269 ( .A1(n26433), .A2(n26434), .A3(n26435), .A4(n26436), .Z(n26432)
         );
  NR4D0 U9270 ( .A1(n26437), .A2(n26438), .A3(n26439), .A4(n26440), .ZN(n26436) );
  OAI222D0 U9271 ( .A1(n24979), .A2(n15585), .B1(n24980), .B2(n4440), .C1(
        n24964), .C2(n2232), .ZN(n26440) );
  OAI222D0 U9272 ( .A1(n24920), .A2(n2520), .B1(n24981), .B2(n5160), .C1(
        n24963), .C2(n2424), .ZN(n26439) );
  OAI222D0 U9273 ( .A1(n24982), .A2(n4920), .B1(n24983), .B2(n4968), .C1(
        n24984), .C2(n4872), .ZN(n26438) );
  OAI222D0 U9274 ( .A1(n24985), .A2(n4392), .B1(n24986), .B2(n3768), .C1(
        n24987), .C2(n4344), .ZN(n26437) );
  NR4D0 U9275 ( .A1(n26441), .A2(n26442), .A3(n26443), .A4(n26444), .ZN(n26435) );
  OAI22D0 U9276 ( .A1(n24922), .A2(n2808), .B1(n24992), .B2(n3720), .ZN(n26444) );
  OAI222D0 U9277 ( .A1(n24993), .A2(n18028), .B1(n24962), .B2(n2760), .C1(
        n24994), .C2(n18029), .ZN(n26443) );
  OAI222D0 U9278 ( .A1(n24995), .A2(n5208), .B1(n24961), .B2(n2664), .C1(
        n24921), .C2(n2712), .ZN(n26442) );
  OAI222D0 U9279 ( .A1(n24927), .A2(n3144), .B1(n24996), .B2(n4776), .C1(
        n24997), .C2(n15584), .ZN(n26441) );
  NR4D0 U9280 ( .A1(n26445), .A2(n26446), .A3(n26447), .A4(n26448), .ZN(n26434) );
  OAI22D0 U9281 ( .A1(n24928), .A2(n3192), .B1(n24926), .B2(n3096), .ZN(n26448) );
  OAI222D0 U9282 ( .A1(n25002), .A2(n3432), .B1(n24929), .B2(n3240), .C1(
        n24933), .C2(n2328), .ZN(n26447) );
  OAI222D0 U9283 ( .A1(n25003), .A2(n3576), .B1(n25004), .B2(n3480), .C1(
        n25005), .C2(n3528), .ZN(n26446) );
  OAI222D0 U9284 ( .A1(n24965), .A2(n2568), .B1(n25006), .B2(n3624), .C1(
        n25007), .C2(n3672), .ZN(n26445) );
  NR4D0 U9285 ( .A1(n26449), .A2(n26450), .A3(n26451), .A4(n26452), .ZN(n26433) );
  OAI22D0 U9286 ( .A1(n25012), .A2(n5112), .B1(n24966), .B2(n2280), .ZN(n26452) );
  OAI222D0 U9287 ( .A1(n24925), .A2(n3048), .B1(n24923), .B2(n2952), .C1(
        n24960), .C2(n2856), .ZN(n26451) );
  OAI222D0 U9288 ( .A1(n25013), .A2(n5496), .B1(n25014), .B2(n5544), .C1(
        n24924), .C2(n3000), .ZN(n26450) );
  OAI222D0 U9289 ( .A1(n25015), .A2(n6072), .B1(n25016), .B2(n5976), .C1(
        n25017), .C2(n6120), .ZN(n26449) );
  INR4D0 U9290 ( .A1(n26453), .B1(n26454), .B2(n26455), .B3(n26456), .ZN(
        n26431) );
  OAI222D0 U9291 ( .A1(n25022), .A2(n5448), .B1(n25023), .B2(n6312), .C1(
        n25024), .C2(n5400), .ZN(n26456) );
  OAI222D0 U9292 ( .A1(n25025), .A2(n4488), .B1(n25026), .B2(n24661), .C1(
        n25027), .C2(n5592), .ZN(n26455) );
  OR4D0 U9293 ( .A1(n26457), .A2(n26458), .A3(n26459), .A4(n26460), .Z(n26454)
         );
  OAI222D0 U9294 ( .A1(n25032), .A2(n4584), .B1(n25033), .B2(n5304), .C1(
        n25034), .C2(n6216), .ZN(n26460) );
  OAI222D0 U9295 ( .A1(n25035), .A2(n6168), .B1(n25036), .B2(n4536), .C1(
        n25037), .C2(n5352), .ZN(n26459) );
  OAI22D0 U9296 ( .A1(n27175), .A2(n25038), .B1(n27174), .B2(n25039), .ZN(
        n26458) );
  OAI222D0 U9297 ( .A1(n24846), .A2(n25040), .B1(n25041), .B2(n5832), .C1(
        n25042), .C2(n5784), .ZN(n26457) );
  CKND0 U9298 ( .I(\Mem[44][34] ), .ZN(n24846) );
  AOI221D0 U9299 ( .A1(n27172), .A2(n25043), .B1(n27173), .B2(n25044), .C(
        n26461), .ZN(n26453) );
  OAI222D0 U9300 ( .A1(n25046), .A2(n6024), .B1(n24847), .B2(n25047), .C1(
        n25048), .C2(n4680), .ZN(n26461) );
  CKND0 U9301 ( .I(\Mem[45][34] ), .ZN(n24847) );
  NR4D0 U9302 ( .A1(n26462), .A2(n26463), .A3(n26464), .A4(n26465), .ZN(n26430) );
  OAI22D0 U9303 ( .A1(n25053), .A2(n5880), .B1(n25054), .B2(n5688), .ZN(n26465) );
  OAI222D0 U9304 ( .A1(n25055), .A2(n3816), .B1(n25056), .B2(n3864), .C1(
        n25057), .C2(n5928), .ZN(n26464) );
  OAI222D0 U9305 ( .A1(n25058), .A2(n3960), .B1(n25059), .B2(n4008), .C1(
        n25060), .C2(n3912), .ZN(n26463) );
  OAI222D0 U9306 ( .A1(n25061), .A2(n4104), .B1(n25062), .B2(n4152), .C1(
        n25063), .C2(n4056), .ZN(n26462) );
  NR4D0 U9307 ( .A1(n26466), .A2(n26467), .A3(n26468), .A4(n26469), .ZN(n26429) );
  OAI22D0 U9308 ( .A1(n25068), .A2(n2376), .B1(n25069), .B2(n2904), .ZN(n26469) );
  OAI222D0 U9309 ( .A1(n25070), .A2(n2472), .B1(n25071), .B2(n4296), .C1(
        n25072), .C2(n2616), .ZN(n26468) );
  OAI222D0 U9310 ( .A1(n25073), .A2(n4248), .B1(n24930), .B2(n3288), .C1(
        n25074), .C2(n4200), .ZN(n26467) );
  OAI222D0 U9311 ( .A1(n24932), .A2(n3384), .B1(n25075), .B2(n4824), .C1(
        n24931), .C2(n3336), .ZN(n26466) );
  ND4D0 U9312 ( .A1(n26470), .A2(n26471), .A3(n26472), .A4(n26473), .ZN(n2182)
         );
  AN4D0 U9313 ( .A1(n26474), .A2(n26475), .A3(n26476), .A4(n26477), .Z(n26473)
         );
  NR4D0 U9314 ( .A1(n26478), .A2(n26479), .A3(n26480), .A4(n26481), .ZN(n26477) );
  OAI222D0 U9315 ( .A1(n24979), .A2(n15589), .B1(n24980), .B2(n4439), .C1(
        n24964), .C2(n2231), .ZN(n26481) );
  OAI222D0 U9316 ( .A1(n24920), .A2(n2519), .B1(n24981), .B2(n5159), .C1(
        n24963), .C2(n2423), .ZN(n26480) );
  OAI222D0 U9317 ( .A1(n24982), .A2(n4919), .B1(n24983), .B2(n4967), .C1(
        n24984), .C2(n4871), .ZN(n26479) );
  OAI222D0 U9318 ( .A1(n24985), .A2(n4391), .B1(n24986), .B2(n3767), .C1(
        n24987), .C2(n4343), .ZN(n26478) );
  NR4D0 U9319 ( .A1(n26482), .A2(n26483), .A3(n26484), .A4(n26485), .ZN(n26476) );
  OAI22D0 U9320 ( .A1(n24922), .A2(n2807), .B1(n24992), .B2(n3719), .ZN(n26485) );
  OAI222D0 U9321 ( .A1(n24993), .A2(n18031), .B1(n24962), .B2(n2759), .C1(
        n24994), .C2(n18032), .ZN(n26484) );
  OAI222D0 U9322 ( .A1(n24995), .A2(n5207), .B1(n24961), .B2(n2663), .C1(
        n24921), .C2(n2711), .ZN(n26483) );
  OAI222D0 U9323 ( .A1(n24927), .A2(n3143), .B1(n24996), .B2(n4775), .C1(
        n24997), .C2(n15588), .ZN(n26482) );
  NR4D0 U9324 ( .A1(n26486), .A2(n26487), .A3(n26488), .A4(n26489), .ZN(n26475) );
  OAI22D0 U9325 ( .A1(n24928), .A2(n3191), .B1(n24926), .B2(n3095), .ZN(n26489) );
  OAI222D0 U9326 ( .A1(n25002), .A2(n3431), .B1(n24929), .B2(n3239), .C1(
        n24933), .C2(n2327), .ZN(n26488) );
  OAI222D0 U9327 ( .A1(n25003), .A2(n3575), .B1(n25004), .B2(n3479), .C1(
        n25005), .C2(n3527), .ZN(n26487) );
  OAI222D0 U9328 ( .A1(n24965), .A2(n2567), .B1(n25006), .B2(n3623), .C1(
        n25007), .C2(n3671), .ZN(n26486) );
  NR4D0 U9329 ( .A1(n26490), .A2(n26491), .A3(n26492), .A4(n26493), .ZN(n26474) );
  OAI22D0 U9330 ( .A1(n25012), .A2(n5111), .B1(n24966), .B2(n2279), .ZN(n26493) );
  OAI222D0 U9331 ( .A1(n24925), .A2(n3047), .B1(n24923), .B2(n2951), .C1(
        n24960), .C2(n2855), .ZN(n26492) );
  OAI222D0 U9332 ( .A1(n25013), .A2(n5495), .B1(n25014), .B2(n5543), .C1(
        n24924), .C2(n2999), .ZN(n26491) );
  OAI222D0 U9333 ( .A1(n25015), .A2(n6071), .B1(n25016), .B2(n5975), .C1(
        n25017), .C2(n6119), .ZN(n26490) );
  INR4D0 U9334 ( .A1(n26494), .B1(n26495), .B2(n26496), .B3(n26497), .ZN(
        n26472) );
  OAI222D0 U9335 ( .A1(n25022), .A2(n5447), .B1(n25023), .B2(n6311), .C1(
        n25024), .C2(n5399), .ZN(n26497) );
  OAI222D0 U9336 ( .A1(n25025), .A2(n4487), .B1(n25026), .B2(n24664), .C1(
        n25027), .C2(n5591), .ZN(n26496) );
  OR4D0 U9337 ( .A1(n26498), .A2(n26499), .A3(n26500), .A4(n26501), .Z(n26495)
         );
  OAI222D0 U9338 ( .A1(n25032), .A2(n4583), .B1(n25033), .B2(n5303), .C1(
        n25034), .C2(n6215), .ZN(n26501) );
  OAI222D0 U9339 ( .A1(n25035), .A2(n6167), .B1(n25036), .B2(n4535), .C1(
        n25037), .C2(n5351), .ZN(n26500) );
  OAI22D0 U9340 ( .A1(n27179), .A2(n25038), .B1(n27178), .B2(n25039), .ZN(
        n26499) );
  OAI222D0 U9341 ( .A1(n24844), .A2(n25040), .B1(n25041), .B2(n5831), .C1(
        n25042), .C2(n5783), .ZN(n26498) );
  CKND0 U9342 ( .I(\Mem[44][35] ), .ZN(n24844) );
  AOI221D0 U9343 ( .A1(n27176), .A2(n25043), .B1(n27177), .B2(n25044), .C(
        n26502), .ZN(n26494) );
  OAI222D0 U9344 ( .A1(n25046), .A2(n6023), .B1(n24845), .B2(n25047), .C1(
        n25048), .C2(n4679), .ZN(n26502) );
  CKND0 U9345 ( .I(\Mem[45][35] ), .ZN(n24845) );
  NR4D0 U9346 ( .A1(n26503), .A2(n26504), .A3(n26505), .A4(n26506), .ZN(n26471) );
  OAI22D0 U9347 ( .A1(n25053), .A2(n5879), .B1(n25054), .B2(n5687), .ZN(n26506) );
  OAI222D0 U9348 ( .A1(n25055), .A2(n3815), .B1(n25056), .B2(n3863), .C1(
        n25057), .C2(n5927), .ZN(n26505) );
  OAI222D0 U9349 ( .A1(n25058), .A2(n3959), .B1(n25059), .B2(n4007), .C1(
        n25060), .C2(n3911), .ZN(n26504) );
  OAI222D0 U9350 ( .A1(n25061), .A2(n4103), .B1(n25062), .B2(n4151), .C1(
        n25063), .C2(n4055), .ZN(n26503) );
  NR4D0 U9351 ( .A1(n26507), .A2(n26508), .A3(n26509), .A4(n26510), .ZN(n26470) );
  OAI22D0 U9352 ( .A1(n25068), .A2(n2375), .B1(n25069), .B2(n2903), .ZN(n26510) );
  OAI222D0 U9353 ( .A1(n25070), .A2(n2471), .B1(n25071), .B2(n4295), .C1(
        n25072), .C2(n2615), .ZN(n26509) );
  OAI222D0 U9354 ( .A1(n25073), .A2(n4247), .B1(n24930), .B2(n3287), .C1(
        n25074), .C2(n4199), .ZN(n26508) );
  OAI222D0 U9355 ( .A1(n24932), .A2(n3383), .B1(n25075), .B2(n4823), .C1(
        n24931), .C2(n3335), .ZN(n26507) );
  ND4D0 U9356 ( .A1(n26511), .A2(n26512), .A3(n26513), .A4(n26514), .ZN(n2181)
         );
  AN4D0 U9357 ( .A1(n26515), .A2(n26516), .A3(n26517), .A4(n26518), .Z(n26514)
         );
  NR4D0 U9358 ( .A1(n26519), .A2(n26520), .A3(n26521), .A4(n26522), .ZN(n26518) );
  OAI222D0 U9359 ( .A1(n24979), .A2(n15593), .B1(n24980), .B2(n4438), .C1(
        n24964), .C2(n2230), .ZN(n26522) );
  OAI222D0 U9360 ( .A1(n24920), .A2(n2518), .B1(n24981), .B2(n5158), .C1(
        n24963), .C2(n2422), .ZN(n26521) );
  OAI222D0 U9361 ( .A1(n24982), .A2(n4918), .B1(n24983), .B2(n4966), .C1(
        n24984), .C2(n4870), .ZN(n26520) );
  OAI222D0 U9362 ( .A1(n24985), .A2(n4390), .B1(n24986), .B2(n3766), .C1(
        n24987), .C2(n4342), .ZN(n26519) );
  NR4D0 U9363 ( .A1(n26523), .A2(n26524), .A3(n26525), .A4(n26526), .ZN(n26517) );
  OAI22D0 U9364 ( .A1(n24922), .A2(n2806), .B1(n24992), .B2(n3718), .ZN(n26526) );
  OAI222D0 U9365 ( .A1(n24993), .A2(n18034), .B1(n24962), .B2(n2758), .C1(
        n24994), .C2(n18035), .ZN(n26525) );
  OAI222D0 U9366 ( .A1(n24995), .A2(n5206), .B1(n24961), .B2(n2662), .C1(
        n24921), .C2(n2710), .ZN(n26524) );
  OAI222D0 U9367 ( .A1(n24927), .A2(n3142), .B1(n24996), .B2(n4774), .C1(
        n24997), .C2(n15592), .ZN(n26523) );
  NR4D0 U9368 ( .A1(n26527), .A2(n26528), .A3(n26529), .A4(n26530), .ZN(n26516) );
  OAI22D0 U9369 ( .A1(n24928), .A2(n3190), .B1(n24926), .B2(n3094), .ZN(n26530) );
  OAI222D0 U9370 ( .A1(n25002), .A2(n3430), .B1(n24929), .B2(n3238), .C1(
        n24933), .C2(n2326), .ZN(n26529) );
  OAI222D0 U9371 ( .A1(n25003), .A2(n3574), .B1(n25004), .B2(n3478), .C1(
        n25005), .C2(n3526), .ZN(n26528) );
  OAI222D0 U9372 ( .A1(n24965), .A2(n2566), .B1(n25006), .B2(n3622), .C1(
        n25007), .C2(n3670), .ZN(n26527) );
  NR4D0 U9373 ( .A1(n26531), .A2(n26532), .A3(n26533), .A4(n26534), .ZN(n26515) );
  OAI22D0 U9374 ( .A1(n25012), .A2(n5110), .B1(n24966), .B2(n2278), .ZN(n26534) );
  OAI222D0 U9375 ( .A1(n24925), .A2(n3046), .B1(n24923), .B2(n2950), .C1(
        n24960), .C2(n2854), .ZN(n26533) );
  OAI222D0 U9376 ( .A1(n25013), .A2(n5494), .B1(n25014), .B2(n5542), .C1(
        n24924), .C2(n2998), .ZN(n26532) );
  OAI222D0 U9377 ( .A1(n25015), .A2(n6070), .B1(n25016), .B2(n5974), .C1(
        n25017), .C2(n6118), .ZN(n26531) );
  INR4D0 U9378 ( .A1(n26535), .B1(n26536), .B2(n26537), .B3(n26538), .ZN(
        n26513) );
  OAI222D0 U9379 ( .A1(n25022), .A2(n5446), .B1(n25023), .B2(n6310), .C1(
        n25024), .C2(n5398), .ZN(n26538) );
  OAI222D0 U9380 ( .A1(n25025), .A2(n4486), .B1(n25026), .B2(n24667), .C1(
        n25027), .C2(n5590), .ZN(n26537) );
  OR4D0 U9381 ( .A1(n26539), .A2(n26540), .A3(n26541), .A4(n26542), .Z(n26536)
         );
  OAI222D0 U9382 ( .A1(n25032), .A2(n4582), .B1(n25033), .B2(n5302), .C1(
        n25034), .C2(n6214), .ZN(n26542) );
  OAI222D0 U9383 ( .A1(n25035), .A2(n6166), .B1(n25036), .B2(n4534), .C1(
        n25037), .C2(n5350), .ZN(n26541) );
  OAI22D0 U9384 ( .A1(n27183), .A2(n25038), .B1(n27182), .B2(n25039), .ZN(
        n26540) );
  OAI222D0 U9385 ( .A1(n24842), .A2(n25040), .B1(n25041), .B2(n5830), .C1(
        n25042), .C2(n5782), .ZN(n26539) );
  CKND0 U9386 ( .I(\Mem[44][36] ), .ZN(n24842) );
  AOI221D0 U9387 ( .A1(n27180), .A2(n25043), .B1(n27181), .B2(n25044), .C(
        n26543), .ZN(n26535) );
  OAI222D0 U9388 ( .A1(n25046), .A2(n6022), .B1(n24843), .B2(n25047), .C1(
        n25048), .C2(n4678), .ZN(n26543) );
  CKND0 U9389 ( .I(\Mem[45][36] ), .ZN(n24843) );
  NR4D0 U9390 ( .A1(n26544), .A2(n26545), .A3(n26546), .A4(n26547), .ZN(n26512) );
  OAI22D0 U9391 ( .A1(n25053), .A2(n5878), .B1(n25054), .B2(n5686), .ZN(n26547) );
  OAI222D0 U9392 ( .A1(n25055), .A2(n3814), .B1(n25056), .B2(n3862), .C1(
        n25057), .C2(n5926), .ZN(n26546) );
  OAI222D0 U9393 ( .A1(n25058), .A2(n3958), .B1(n25059), .B2(n4006), .C1(
        n25060), .C2(n3910), .ZN(n26545) );
  OAI222D0 U9394 ( .A1(n25061), .A2(n4102), .B1(n25062), .B2(n4150), .C1(
        n25063), .C2(n4054), .ZN(n26544) );
  NR4D0 U9395 ( .A1(n26548), .A2(n26549), .A3(n26550), .A4(n26551), .ZN(n26511) );
  OAI22D0 U9396 ( .A1(n25068), .A2(n2374), .B1(n25069), .B2(n2902), .ZN(n26551) );
  OAI222D0 U9397 ( .A1(n25070), .A2(n2470), .B1(n25071), .B2(n4294), .C1(
        n25072), .C2(n2614), .ZN(n26550) );
  OAI222D0 U9398 ( .A1(n25073), .A2(n4246), .B1(n24930), .B2(n3286), .C1(
        n25074), .C2(n4198), .ZN(n26549) );
  OAI222D0 U9399 ( .A1(n24932), .A2(n3382), .B1(n25075), .B2(n4822), .C1(
        n24931), .C2(n3334), .ZN(n26548) );
  ND4D0 U9400 ( .A1(n26552), .A2(n26553), .A3(n26554), .A4(n26555), .ZN(n2180)
         );
  AN4D0 U9401 ( .A1(n26556), .A2(n26557), .A3(n26558), .A4(n26559), .Z(n26555)
         );
  NR4D0 U9402 ( .A1(n26560), .A2(n26561), .A3(n26562), .A4(n26563), .ZN(n26559) );
  OAI222D0 U9403 ( .A1(n24979), .A2(n15597), .B1(n24980), .B2(n4437), .C1(
        n24964), .C2(n2229), .ZN(n26563) );
  OAI222D0 U9404 ( .A1(n24920), .A2(n2517), .B1(n24981), .B2(n5157), .C1(
        n24963), .C2(n2421), .ZN(n26562) );
  OAI222D0 U9405 ( .A1(n24982), .A2(n4917), .B1(n24983), .B2(n4965), .C1(
        n24984), .C2(n4869), .ZN(n26561) );
  OAI222D0 U9406 ( .A1(n24985), .A2(n4389), .B1(n24986), .B2(n3765), .C1(
        n24987), .C2(n4341), .ZN(n26560) );
  NR4D0 U9407 ( .A1(n26564), .A2(n26565), .A3(n26566), .A4(n26567), .ZN(n26558) );
  OAI22D0 U9408 ( .A1(n24922), .A2(n2805), .B1(n24992), .B2(n3717), .ZN(n26567) );
  OAI222D0 U9409 ( .A1(n24993), .A2(n18037), .B1(n24962), .B2(n2757), .C1(
        n24994), .C2(n18038), .ZN(n26566) );
  OAI222D0 U9410 ( .A1(n24995), .A2(n5205), .B1(n24961), .B2(n2661), .C1(
        n24921), .C2(n2709), .ZN(n26565) );
  OAI222D0 U9411 ( .A1(n24927), .A2(n3141), .B1(n24996), .B2(n4773), .C1(
        n24997), .C2(n15596), .ZN(n26564) );
  NR4D0 U9412 ( .A1(n26568), .A2(n26569), .A3(n26570), .A4(n26571), .ZN(n26557) );
  OAI22D0 U9413 ( .A1(n24928), .A2(n3189), .B1(n24926), .B2(n3093), .ZN(n26571) );
  OAI222D0 U9414 ( .A1(n25002), .A2(n3429), .B1(n24929), .B2(n3237), .C1(
        n24933), .C2(n2325), .ZN(n26570) );
  OAI222D0 U9415 ( .A1(n25003), .A2(n3573), .B1(n25004), .B2(n3477), .C1(
        n25005), .C2(n3525), .ZN(n26569) );
  OAI222D0 U9416 ( .A1(n24965), .A2(n2565), .B1(n25006), .B2(n3621), .C1(
        n25007), .C2(n3669), .ZN(n26568) );
  NR4D0 U9417 ( .A1(n26572), .A2(n26573), .A3(n26574), .A4(n26575), .ZN(n26556) );
  OAI22D0 U9418 ( .A1(n25012), .A2(n5109), .B1(n24966), .B2(n2277), .ZN(n26575) );
  OAI222D0 U9419 ( .A1(n24925), .A2(n3045), .B1(n24923), .B2(n2949), .C1(
        n24960), .C2(n2853), .ZN(n26574) );
  OAI222D0 U9420 ( .A1(n25013), .A2(n5493), .B1(n25014), .B2(n5541), .C1(
        n24924), .C2(n2997), .ZN(n26573) );
  OAI222D0 U9421 ( .A1(n25015), .A2(n6069), .B1(n25016), .B2(n5973), .C1(
        n25017), .C2(n6117), .ZN(n26572) );
  INR4D0 U9422 ( .A1(n26576), .B1(n26577), .B2(n26578), .B3(n26579), .ZN(
        n26554) );
  OAI222D0 U9423 ( .A1(n25022), .A2(n5445), .B1(n25023), .B2(n6309), .C1(
        n25024), .C2(n5397), .ZN(n26579) );
  OAI222D0 U9424 ( .A1(n25025), .A2(n4485), .B1(n25026), .B2(n24670), .C1(
        n25027), .C2(n5589), .ZN(n26578) );
  OR4D0 U9425 ( .A1(n26580), .A2(n26581), .A3(n26582), .A4(n26583), .Z(n26577)
         );
  OAI222D0 U9426 ( .A1(n25032), .A2(n4581), .B1(n25033), .B2(n5301), .C1(
        n25034), .C2(n6213), .ZN(n26583) );
  OAI222D0 U9427 ( .A1(n25035), .A2(n6165), .B1(n25036), .B2(n4533), .C1(
        n25037), .C2(n5349), .ZN(n26582) );
  OAI22D0 U9428 ( .A1(n27187), .A2(n25038), .B1(n27186), .B2(n25039), .ZN(
        n26581) );
  OAI222D0 U9429 ( .A1(n24840), .A2(n25040), .B1(n25041), .B2(n5829), .C1(
        n25042), .C2(n5781), .ZN(n26580) );
  CKND0 U9430 ( .I(\Mem[44][37] ), .ZN(n24840) );
  AOI221D0 U9431 ( .A1(n27184), .A2(n25043), .B1(n27185), .B2(n25044), .C(
        n26584), .ZN(n26576) );
  OAI222D0 U9432 ( .A1(n25046), .A2(n6021), .B1(n24841), .B2(n25047), .C1(
        n25048), .C2(n4677), .ZN(n26584) );
  CKND0 U9433 ( .I(\Mem[45][37] ), .ZN(n24841) );
  NR4D0 U9434 ( .A1(n26585), .A2(n26586), .A3(n26587), .A4(n26588), .ZN(n26553) );
  OAI22D0 U9435 ( .A1(n25053), .A2(n5877), .B1(n25054), .B2(n5685), .ZN(n26588) );
  OAI222D0 U9436 ( .A1(n25055), .A2(n3813), .B1(n25056), .B2(n3861), .C1(
        n25057), .C2(n5925), .ZN(n26587) );
  OAI222D0 U9437 ( .A1(n25058), .A2(n3957), .B1(n25059), .B2(n4005), .C1(
        n25060), .C2(n3909), .ZN(n26586) );
  OAI222D0 U9438 ( .A1(n25061), .A2(n4101), .B1(n25062), .B2(n4149), .C1(
        n25063), .C2(n4053), .ZN(n26585) );
  NR4D0 U9439 ( .A1(n26589), .A2(n26590), .A3(n26591), .A4(n26592), .ZN(n26552) );
  OAI22D0 U9440 ( .A1(n25068), .A2(n2373), .B1(n25069), .B2(n2901), .ZN(n26592) );
  OAI222D0 U9441 ( .A1(n25070), .A2(n2469), .B1(n25071), .B2(n4293), .C1(
        n25072), .C2(n2613), .ZN(n26591) );
  OAI222D0 U9442 ( .A1(n25073), .A2(n4245), .B1(n24930), .B2(n3285), .C1(
        n25074), .C2(n4197), .ZN(n26590) );
  OAI222D0 U9443 ( .A1(n24932), .A2(n3381), .B1(n25075), .B2(n4821), .C1(
        n24931), .C2(n3333), .ZN(n26589) );
  ND4D0 U9444 ( .A1(n26593), .A2(n26594), .A3(n26595), .A4(n26596), .ZN(n2179)
         );
  AN4D0 U9445 ( .A1(n26597), .A2(n26598), .A3(n26599), .A4(n26600), .Z(n26596)
         );
  NR4D0 U9446 ( .A1(n26601), .A2(n26602), .A3(n26603), .A4(n26604), .ZN(n26600) );
  OAI222D0 U9447 ( .A1(n24979), .A2(n15601), .B1(n24980), .B2(n4436), .C1(
        n24964), .C2(n2228), .ZN(n26604) );
  OAI222D0 U9448 ( .A1(n24920), .A2(n2516), .B1(n24981), .B2(n5156), .C1(
        n24963), .C2(n2420), .ZN(n26603) );
  OAI222D0 U9449 ( .A1(n24982), .A2(n4916), .B1(n24983), .B2(n4964), .C1(
        n24984), .C2(n4868), .ZN(n26602) );
  OAI222D0 U9450 ( .A1(n24985), .A2(n4388), .B1(n24986), .B2(n3764), .C1(
        n24987), .C2(n4340), .ZN(n26601) );
  NR4D0 U9451 ( .A1(n26605), .A2(n26606), .A3(n26607), .A4(n26608), .ZN(n26599) );
  OAI22D0 U9452 ( .A1(n24922), .A2(n2804), .B1(n24992), .B2(n3716), .ZN(n26608) );
  OAI222D0 U9453 ( .A1(n24993), .A2(n18040), .B1(n24962), .B2(n2756), .C1(
        n24994), .C2(n18041), .ZN(n26607) );
  OAI222D0 U9454 ( .A1(n24995), .A2(n5204), .B1(n24961), .B2(n2660), .C1(
        n24921), .C2(n2708), .ZN(n26606) );
  OAI222D0 U9455 ( .A1(n24927), .A2(n3140), .B1(n24996), .B2(n4772), .C1(
        n24997), .C2(n15600), .ZN(n26605) );
  NR4D0 U9456 ( .A1(n26609), .A2(n26610), .A3(n26611), .A4(n26612), .ZN(n26598) );
  OAI22D0 U9457 ( .A1(n24928), .A2(n3188), .B1(n24926), .B2(n3092), .ZN(n26612) );
  OAI222D0 U9458 ( .A1(n25002), .A2(n3428), .B1(n24929), .B2(n3236), .C1(
        n24933), .C2(n2324), .ZN(n26611) );
  OAI222D0 U9459 ( .A1(n25003), .A2(n3572), .B1(n25004), .B2(n3476), .C1(
        n25005), .C2(n3524), .ZN(n26610) );
  OAI222D0 U9460 ( .A1(n24965), .A2(n2564), .B1(n25006), .B2(n3620), .C1(
        n25007), .C2(n3668), .ZN(n26609) );
  NR4D0 U9461 ( .A1(n26613), .A2(n26614), .A3(n26615), .A4(n26616), .ZN(n26597) );
  OAI22D0 U9462 ( .A1(n25012), .A2(n5108), .B1(n24966), .B2(n2276), .ZN(n26616) );
  OAI222D0 U9463 ( .A1(n24925), .A2(n3044), .B1(n24923), .B2(n2948), .C1(
        n24960), .C2(n2852), .ZN(n26615) );
  OAI222D0 U9464 ( .A1(n25013), .A2(n5492), .B1(n25014), .B2(n5540), .C1(
        n24924), .C2(n2996), .ZN(n26614) );
  OAI222D0 U9465 ( .A1(n25015), .A2(n6068), .B1(n25016), .B2(n5972), .C1(
        n25017), .C2(n6116), .ZN(n26613) );
  INR4D0 U9466 ( .A1(n26617), .B1(n26618), .B2(n26619), .B3(n26620), .ZN(
        n26595) );
  OAI222D0 U9467 ( .A1(n25022), .A2(n5444), .B1(n25023), .B2(n6308), .C1(
        n25024), .C2(n5396), .ZN(n26620) );
  OAI222D0 U9468 ( .A1(n25025), .A2(n4484), .B1(n25026), .B2(n24673), .C1(
        n25027), .C2(n5588), .ZN(n26619) );
  OR4D0 U9469 ( .A1(n26621), .A2(n26622), .A3(n26623), .A4(n26624), .Z(n26618)
         );
  OAI222D0 U9470 ( .A1(n25032), .A2(n4580), .B1(n25033), .B2(n5300), .C1(
        n25034), .C2(n6212), .ZN(n26624) );
  OAI222D0 U9471 ( .A1(n25035), .A2(n6164), .B1(n25036), .B2(n4532), .C1(
        n25037), .C2(n5348), .ZN(n26623) );
  OAI22D0 U9472 ( .A1(n27191), .A2(n25038), .B1(n27190), .B2(n25039), .ZN(
        n26622) );
  OAI222D0 U9473 ( .A1(n24838), .A2(n25040), .B1(n25041), .B2(n5828), .C1(
        n25042), .C2(n5780), .ZN(n26621) );
  CKND0 U9474 ( .I(\Mem[44][38] ), .ZN(n24838) );
  AOI221D0 U9475 ( .A1(n27188), .A2(n25043), .B1(n27189), .B2(n25044), .C(
        n26625), .ZN(n26617) );
  OAI222D0 U9476 ( .A1(n25046), .A2(n6020), .B1(n24839), .B2(n25047), .C1(
        n25048), .C2(n4676), .ZN(n26625) );
  CKND0 U9477 ( .I(\Mem[45][38] ), .ZN(n24839) );
  NR4D0 U9478 ( .A1(n26626), .A2(n26627), .A3(n26628), .A4(n26629), .ZN(n26594) );
  OAI22D0 U9479 ( .A1(n25053), .A2(n5876), .B1(n25054), .B2(n5684), .ZN(n26629) );
  OAI222D0 U9480 ( .A1(n25055), .A2(n3812), .B1(n25056), .B2(n3860), .C1(
        n25057), .C2(n5924), .ZN(n26628) );
  OAI222D0 U9481 ( .A1(n25058), .A2(n3956), .B1(n25059), .B2(n4004), .C1(
        n25060), .C2(n3908), .ZN(n26627) );
  OAI222D0 U9482 ( .A1(n25061), .A2(n4100), .B1(n25062), .B2(n4148), .C1(
        n25063), .C2(n4052), .ZN(n26626) );
  NR4D0 U9483 ( .A1(n26630), .A2(n26631), .A3(n26632), .A4(n26633), .ZN(n26593) );
  OAI22D0 U9484 ( .A1(n25068), .A2(n2372), .B1(n25069), .B2(n2900), .ZN(n26633) );
  OAI222D0 U9485 ( .A1(n25070), .A2(n2468), .B1(n25071), .B2(n4292), .C1(
        n25072), .C2(n2612), .ZN(n26632) );
  OAI222D0 U9486 ( .A1(n25073), .A2(n4244), .B1(n24930), .B2(n3284), .C1(
        n25074), .C2(n4196), .ZN(n26631) );
  OAI222D0 U9487 ( .A1(n24932), .A2(n3380), .B1(n25075), .B2(n4820), .C1(
        n24931), .C2(n3332), .ZN(n26630) );
  ND4D0 U9488 ( .A1(n26634), .A2(n26635), .A3(n26636), .A4(n26637), .ZN(n2178)
         );
  AN4D0 U9489 ( .A1(n26638), .A2(n26639), .A3(n26640), .A4(n26641), .Z(n26637)
         );
  NR4D0 U9490 ( .A1(n26642), .A2(n26643), .A3(n26644), .A4(n26645), .ZN(n26641) );
  OAI222D0 U9491 ( .A1(n24979), .A2(n15605), .B1(n24980), .B2(n4435), .C1(
        n24964), .C2(n2227), .ZN(n26645) );
  OAI222D0 U9492 ( .A1(n24920), .A2(n2515), .B1(n24981), .B2(n5155), .C1(
        n24963), .C2(n2419), .ZN(n26644) );
  OAI222D0 U9493 ( .A1(n24982), .A2(n4915), .B1(n24983), .B2(n4963), .C1(
        n24984), .C2(n4867), .ZN(n26643) );
  OAI222D0 U9494 ( .A1(n24985), .A2(n4387), .B1(n24986), .B2(n3763), .C1(
        n24987), .C2(n4339), .ZN(n26642) );
  NR4D0 U9495 ( .A1(n26646), .A2(n26647), .A3(n26648), .A4(n26649), .ZN(n26640) );
  OAI22D0 U9496 ( .A1(n24922), .A2(n2803), .B1(n24992), .B2(n3715), .ZN(n26649) );
  OAI222D0 U9497 ( .A1(n24993), .A2(n18043), .B1(n24962), .B2(n2755), .C1(
        n24994), .C2(n18044), .ZN(n26648) );
  OAI222D0 U9498 ( .A1(n24995), .A2(n5203), .B1(n24961), .B2(n2659), .C1(
        n24921), .C2(n2707), .ZN(n26647) );
  OAI222D0 U9499 ( .A1(n24927), .A2(n3139), .B1(n24996), .B2(n4771), .C1(
        n24997), .C2(n15604), .ZN(n26646) );
  NR4D0 U9500 ( .A1(n26650), .A2(n26651), .A3(n26652), .A4(n26653), .ZN(n26639) );
  OAI22D0 U9501 ( .A1(n24928), .A2(n3187), .B1(n24926), .B2(n3091), .ZN(n26653) );
  OAI222D0 U9502 ( .A1(n25002), .A2(n3427), .B1(n24929), .B2(n3235), .C1(
        n24933), .C2(n2323), .ZN(n26652) );
  OAI222D0 U9503 ( .A1(n25003), .A2(n3571), .B1(n25004), .B2(n3475), .C1(
        n25005), .C2(n3523), .ZN(n26651) );
  OAI222D0 U9504 ( .A1(n24965), .A2(n2563), .B1(n25006), .B2(n3619), .C1(
        n25007), .C2(n3667), .ZN(n26650) );
  NR4D0 U9505 ( .A1(n26654), .A2(n26655), .A3(n26656), .A4(n26657), .ZN(n26638) );
  OAI22D0 U9506 ( .A1(n25012), .A2(n5107), .B1(n24966), .B2(n2275), .ZN(n26657) );
  OAI222D0 U9507 ( .A1(n24925), .A2(n3043), .B1(n24923), .B2(n2947), .C1(
        n24960), .C2(n2851), .ZN(n26656) );
  OAI222D0 U9508 ( .A1(n25013), .A2(n5491), .B1(n25014), .B2(n5539), .C1(
        n24924), .C2(n2995), .ZN(n26655) );
  OAI222D0 U9509 ( .A1(n25015), .A2(n6067), .B1(n25016), .B2(n5971), .C1(
        n25017), .C2(n6115), .ZN(n26654) );
  INR4D0 U9510 ( .A1(n26658), .B1(n26659), .B2(n26660), .B3(n26661), .ZN(
        n26636) );
  OAI222D0 U9511 ( .A1(n25022), .A2(n5443), .B1(n25023), .B2(n6307), .C1(
        n25024), .C2(n5395), .ZN(n26661) );
  OAI222D0 U9512 ( .A1(n25025), .A2(n4483), .B1(n25026), .B2(n24676), .C1(
        n25027), .C2(n5587), .ZN(n26660) );
  OR4D0 U9513 ( .A1(n26662), .A2(n26663), .A3(n26664), .A4(n26665), .Z(n26659)
         );
  OAI222D0 U9514 ( .A1(n25032), .A2(n4579), .B1(n25033), .B2(n5299), .C1(
        n25034), .C2(n6211), .ZN(n26665) );
  OAI222D0 U9515 ( .A1(n25035), .A2(n6163), .B1(n25036), .B2(n4531), .C1(
        n25037), .C2(n5347), .ZN(n26664) );
  OAI22D0 U9516 ( .A1(n27195), .A2(n25038), .B1(n27194), .B2(n25039), .ZN(
        n26663) );
  OAI222D0 U9517 ( .A1(n24836), .A2(n25040), .B1(n25041), .B2(n5827), .C1(
        n25042), .C2(n5779), .ZN(n26662) );
  CKND0 U9518 ( .I(\Mem[44][39] ), .ZN(n24836) );
  AOI221D0 U9519 ( .A1(n27192), .A2(n25043), .B1(n27193), .B2(n25044), .C(
        n26666), .ZN(n26658) );
  OAI222D0 U9520 ( .A1(n25046), .A2(n6019), .B1(n24837), .B2(n25047), .C1(
        n25048), .C2(n4675), .ZN(n26666) );
  CKND0 U9521 ( .I(\Mem[45][39] ), .ZN(n24837) );
  NR4D0 U9522 ( .A1(n26667), .A2(n26668), .A3(n26669), .A4(n26670), .ZN(n26635) );
  OAI22D0 U9523 ( .A1(n25053), .A2(n5875), .B1(n25054), .B2(n5683), .ZN(n26670) );
  OAI222D0 U9524 ( .A1(n25055), .A2(n3811), .B1(n25056), .B2(n3859), .C1(
        n25057), .C2(n5923), .ZN(n26669) );
  OAI222D0 U9525 ( .A1(n25058), .A2(n3955), .B1(n25059), .B2(n4003), .C1(
        n25060), .C2(n3907), .ZN(n26668) );
  OAI222D0 U9526 ( .A1(n25061), .A2(n4099), .B1(n25062), .B2(n4147), .C1(
        n25063), .C2(n4051), .ZN(n26667) );
  NR4D0 U9527 ( .A1(n26671), .A2(n26672), .A3(n26673), .A4(n26674), .ZN(n26634) );
  OAI22D0 U9528 ( .A1(n25068), .A2(n2371), .B1(n25069), .B2(n2899), .ZN(n26674) );
  OAI222D0 U9529 ( .A1(n25070), .A2(n2467), .B1(n25071), .B2(n4291), .C1(
        n25072), .C2(n2611), .ZN(n26673) );
  OAI222D0 U9530 ( .A1(n25073), .A2(n4243), .B1(n24930), .B2(n3283), .C1(
        n25074), .C2(n4195), .ZN(n26672) );
  OAI222D0 U9531 ( .A1(n24932), .A2(n3379), .B1(n25075), .B2(n4819), .C1(
        n24931), .C2(n3331), .ZN(n26671) );
  ND4D0 U9532 ( .A1(n26675), .A2(n26676), .A3(n26677), .A4(n26678), .ZN(n2177)
         );
  AN4D0 U9533 ( .A1(n26679), .A2(n26680), .A3(n26681), .A4(n26682), .Z(n26678)
         );
  NR4D0 U9534 ( .A1(n26683), .A2(n26684), .A3(n26685), .A4(n26686), .ZN(n26682) );
  OAI222D0 U9535 ( .A1(n24979), .A2(n15609), .B1(n24980), .B2(n4434), .C1(
        n24964), .C2(n2226), .ZN(n26686) );
  OAI222D0 U9536 ( .A1(n24920), .A2(n2514), .B1(n24981), .B2(n5154), .C1(
        n24963), .C2(n2418), .ZN(n26685) );
  OAI222D0 U9537 ( .A1(n24982), .A2(n4914), .B1(n24983), .B2(n4962), .C1(
        n24984), .C2(n4866), .ZN(n26684) );
  OAI222D0 U9538 ( .A1(n24985), .A2(n4386), .B1(n24986), .B2(n3762), .C1(
        n24987), .C2(n4338), .ZN(n26683) );
  NR4D0 U9539 ( .A1(n26687), .A2(n26688), .A3(n26689), .A4(n26690), .ZN(n26681) );
  OAI22D0 U9540 ( .A1(n24922), .A2(n2802), .B1(n24992), .B2(n3714), .ZN(n26690) );
  OAI222D0 U9541 ( .A1(n24993), .A2(n18046), .B1(n24962), .B2(n2754), .C1(
        n24994), .C2(n18047), .ZN(n26689) );
  OAI222D0 U9542 ( .A1(n24995), .A2(n5202), .B1(n24961), .B2(n2658), .C1(
        n24921), .C2(n2706), .ZN(n26688) );
  OAI222D0 U9543 ( .A1(n24927), .A2(n3138), .B1(n24996), .B2(n4770), .C1(
        n24997), .C2(n15608), .ZN(n26687) );
  NR4D0 U9544 ( .A1(n26691), .A2(n26692), .A3(n26693), .A4(n26694), .ZN(n26680) );
  OAI22D0 U9545 ( .A1(n24928), .A2(n3186), .B1(n24926), .B2(n3090), .ZN(n26694) );
  OAI222D0 U9546 ( .A1(n25002), .A2(n3426), .B1(n24929), .B2(n3234), .C1(
        n24933), .C2(n2322), .ZN(n26693) );
  OAI222D0 U9547 ( .A1(n25003), .A2(n3570), .B1(n25004), .B2(n3474), .C1(
        n25005), .C2(n3522), .ZN(n26692) );
  OAI222D0 U9548 ( .A1(n24965), .A2(n2562), .B1(n25006), .B2(n3618), .C1(
        n25007), .C2(n3666), .ZN(n26691) );
  NR4D0 U9549 ( .A1(n26695), .A2(n26696), .A3(n26697), .A4(n26698), .ZN(n26679) );
  OAI22D0 U9550 ( .A1(n25012), .A2(n5106), .B1(n24966), .B2(n2274), .ZN(n26698) );
  OAI222D0 U9551 ( .A1(n24925), .A2(n3042), .B1(n24923), .B2(n2946), .C1(
        n24960), .C2(n2850), .ZN(n26697) );
  OAI222D0 U9552 ( .A1(n25013), .A2(n5490), .B1(n25014), .B2(n5538), .C1(
        n24924), .C2(n2994), .ZN(n26696) );
  OAI222D0 U9553 ( .A1(n25015), .A2(n6066), .B1(n25016), .B2(n5970), .C1(
        n25017), .C2(n6114), .ZN(n26695) );
  INR4D0 U9554 ( .A1(n26699), .B1(n26700), .B2(n26701), .B3(n26702), .ZN(
        n26677) );
  OAI222D0 U9555 ( .A1(n25022), .A2(n5442), .B1(n25023), .B2(n6306), .C1(
        n25024), .C2(n5394), .ZN(n26702) );
  OAI222D0 U9556 ( .A1(n25025), .A2(n4482), .B1(n25026), .B2(n24679), .C1(
        n25027), .C2(n5586), .ZN(n26701) );
  OR4D0 U9557 ( .A1(n26703), .A2(n26704), .A3(n26705), .A4(n26706), .Z(n26700)
         );
  OAI222D0 U9558 ( .A1(n25032), .A2(n4578), .B1(n25033), .B2(n5298), .C1(
        n25034), .C2(n6210), .ZN(n26706) );
  OAI222D0 U9559 ( .A1(n25035), .A2(n6162), .B1(n25036), .B2(n4530), .C1(
        n25037), .C2(n5346), .ZN(n26705) );
  OAI22D0 U9560 ( .A1(n27199), .A2(n25038), .B1(n27198), .B2(n25039), .ZN(
        n26704) );
  OAI222D0 U9561 ( .A1(n24834), .A2(n25040), .B1(n25041), .B2(n5826), .C1(
        n25042), .C2(n5778), .ZN(n26703) );
  CKND0 U9562 ( .I(\Mem[44][40] ), .ZN(n24834) );
  AOI221D0 U9563 ( .A1(n27196), .A2(n25043), .B1(n27197), .B2(n25044), .C(
        n26707), .ZN(n26699) );
  OAI222D0 U9564 ( .A1(n25046), .A2(n6018), .B1(n24835), .B2(n25047), .C1(
        n25048), .C2(n4674), .ZN(n26707) );
  CKND0 U9565 ( .I(\Mem[45][40] ), .ZN(n24835) );
  NR4D0 U9566 ( .A1(n26708), .A2(n26709), .A3(n26710), .A4(n26711), .ZN(n26676) );
  OAI22D0 U9567 ( .A1(n25053), .A2(n5874), .B1(n25054), .B2(n5682), .ZN(n26711) );
  OAI222D0 U9568 ( .A1(n25055), .A2(n3810), .B1(n25056), .B2(n3858), .C1(
        n25057), .C2(n5922), .ZN(n26710) );
  OAI222D0 U9569 ( .A1(n25058), .A2(n3954), .B1(n25059), .B2(n4002), .C1(
        n25060), .C2(n3906), .ZN(n26709) );
  OAI222D0 U9570 ( .A1(n25061), .A2(n4098), .B1(n25062), .B2(n4146), .C1(
        n25063), .C2(n4050), .ZN(n26708) );
  NR4D0 U9571 ( .A1(n26712), .A2(n26713), .A3(n26714), .A4(n26715), .ZN(n26675) );
  OAI22D0 U9572 ( .A1(n25068), .A2(n2370), .B1(n25069), .B2(n2898), .ZN(n26715) );
  OAI222D0 U9573 ( .A1(n25070), .A2(n2466), .B1(n25071), .B2(n4290), .C1(
        n25072), .C2(n2610), .ZN(n26714) );
  OAI222D0 U9574 ( .A1(n25073), .A2(n4242), .B1(n24930), .B2(n3282), .C1(
        n25074), .C2(n4194), .ZN(n26713) );
  OAI222D0 U9575 ( .A1(n24932), .A2(n3378), .B1(n25075), .B2(n4818), .C1(
        n24931), .C2(n3330), .ZN(n26712) );
  ND4D0 U9576 ( .A1(n26716), .A2(n26717), .A3(n26718), .A4(n26719), .ZN(n2176)
         );
  AN4D0 U9577 ( .A1(n26720), .A2(n26721), .A3(n26722), .A4(n26723), .Z(n26719)
         );
  NR4D0 U9578 ( .A1(n26724), .A2(n26725), .A3(n26726), .A4(n26727), .ZN(n26723) );
  OAI222D0 U9579 ( .A1(n24979), .A2(n15613), .B1(n24980), .B2(n4433), .C1(
        n24964), .C2(n2225), .ZN(n26727) );
  OAI222D0 U9580 ( .A1(n24920), .A2(n2513), .B1(n24981), .B2(n5153), .C1(
        n24963), .C2(n2417), .ZN(n26726) );
  OAI222D0 U9581 ( .A1(n24982), .A2(n4913), .B1(n24983), .B2(n4961), .C1(
        n24984), .C2(n4865), .ZN(n26725) );
  OAI222D0 U9582 ( .A1(n24985), .A2(n4385), .B1(n24986), .B2(n3761), .C1(
        n24987), .C2(n4337), .ZN(n26724) );
  NR4D0 U9583 ( .A1(n26728), .A2(n26729), .A3(n26730), .A4(n26731), .ZN(n26722) );
  OAI22D0 U9584 ( .A1(n24922), .A2(n2801), .B1(n24992), .B2(n3713), .ZN(n26731) );
  OAI222D0 U9585 ( .A1(n24993), .A2(n18049), .B1(n24962), .B2(n2753), .C1(
        n24994), .C2(n18050), .ZN(n26730) );
  OAI222D0 U9586 ( .A1(n24995), .A2(n5201), .B1(n24961), .B2(n2657), .C1(
        n24921), .C2(n2705), .ZN(n26729) );
  OAI222D0 U9587 ( .A1(n24927), .A2(n3137), .B1(n24996), .B2(n4769), .C1(
        n24997), .C2(n15612), .ZN(n26728) );
  NR4D0 U9588 ( .A1(n26732), .A2(n26733), .A3(n26734), .A4(n26735), .ZN(n26721) );
  OAI22D0 U9589 ( .A1(n24928), .A2(n3185), .B1(n24926), .B2(n3089), .ZN(n26735) );
  OAI222D0 U9590 ( .A1(n25002), .A2(n3425), .B1(n24929), .B2(n3233), .C1(
        n24933), .C2(n2321), .ZN(n26734) );
  OAI222D0 U9591 ( .A1(n25003), .A2(n3569), .B1(n25004), .B2(n3473), .C1(
        n25005), .C2(n3521), .ZN(n26733) );
  OAI222D0 U9592 ( .A1(n24965), .A2(n2561), .B1(n25006), .B2(n3617), .C1(
        n25007), .C2(n3665), .ZN(n26732) );
  NR4D0 U9593 ( .A1(n26736), .A2(n26737), .A3(n26738), .A4(n26739), .ZN(n26720) );
  OAI22D0 U9594 ( .A1(n25012), .A2(n5105), .B1(n24966), .B2(n2273), .ZN(n26739) );
  OAI222D0 U9595 ( .A1(n24925), .A2(n3041), .B1(n24923), .B2(n2945), .C1(
        n24960), .C2(n2849), .ZN(n26738) );
  OAI222D0 U9596 ( .A1(n25013), .A2(n5489), .B1(n25014), .B2(n5537), .C1(
        n24924), .C2(n2993), .ZN(n26737) );
  OAI222D0 U9597 ( .A1(n25015), .A2(n6065), .B1(n25016), .B2(n5969), .C1(
        n25017), .C2(n6113), .ZN(n26736) );
  INR4D0 U9598 ( .A1(n26740), .B1(n26741), .B2(n26742), .B3(n26743), .ZN(
        n26718) );
  OAI222D0 U9599 ( .A1(n25022), .A2(n5441), .B1(n25023), .B2(n6305), .C1(
        n25024), .C2(n5393), .ZN(n26743) );
  OAI222D0 U9600 ( .A1(n25025), .A2(n4481), .B1(n25026), .B2(n24682), .C1(
        n25027), .C2(n5585), .ZN(n26742) );
  OR4D0 U9601 ( .A1(n26744), .A2(n26745), .A3(n26746), .A4(n26747), .Z(n26741)
         );
  OAI222D0 U9602 ( .A1(n25032), .A2(n4577), .B1(n25033), .B2(n5297), .C1(
        n25034), .C2(n6209), .ZN(n26747) );
  OAI222D0 U9603 ( .A1(n25035), .A2(n6161), .B1(n25036), .B2(n4529), .C1(
        n25037), .C2(n5345), .ZN(n26746) );
  OAI22D0 U9604 ( .A1(n27203), .A2(n25038), .B1(n27202), .B2(n25039), .ZN(
        n26745) );
  OAI222D0 U9605 ( .A1(n24832), .A2(n25040), .B1(n25041), .B2(n5825), .C1(
        n25042), .C2(n5777), .ZN(n26744) );
  CKND0 U9606 ( .I(\Mem[44][41] ), .ZN(n24832) );
  AOI221D0 U9607 ( .A1(n27200), .A2(n25043), .B1(n27201), .B2(n25044), .C(
        n26748), .ZN(n26740) );
  OAI222D0 U9608 ( .A1(n25046), .A2(n6017), .B1(n24833), .B2(n25047), .C1(
        n25048), .C2(n4673), .ZN(n26748) );
  CKND0 U9609 ( .I(\Mem[45][41] ), .ZN(n24833) );
  NR4D0 U9610 ( .A1(n26749), .A2(n26750), .A3(n26751), .A4(n26752), .ZN(n26717) );
  OAI22D0 U9611 ( .A1(n25053), .A2(n5873), .B1(n25054), .B2(n5681), .ZN(n26752) );
  OAI222D0 U9612 ( .A1(n25055), .A2(n3809), .B1(n25056), .B2(n3857), .C1(
        n25057), .C2(n5921), .ZN(n26751) );
  OAI222D0 U9613 ( .A1(n25058), .A2(n3953), .B1(n25059), .B2(n4001), .C1(
        n25060), .C2(n3905), .ZN(n26750) );
  OAI222D0 U9614 ( .A1(n25061), .A2(n4097), .B1(n25062), .B2(n4145), .C1(
        n25063), .C2(n4049), .ZN(n26749) );
  NR4D0 U9615 ( .A1(n26753), .A2(n26754), .A3(n26755), .A4(n26756), .ZN(n26716) );
  OAI22D0 U9616 ( .A1(n25068), .A2(n2369), .B1(n25069), .B2(n2897), .ZN(n26756) );
  OAI222D0 U9617 ( .A1(n25070), .A2(n2465), .B1(n25071), .B2(n4289), .C1(
        n25072), .C2(n2609), .ZN(n26755) );
  OAI222D0 U9618 ( .A1(n25073), .A2(n4241), .B1(n24930), .B2(n3281), .C1(
        n25074), .C2(n4193), .ZN(n26754) );
  OAI222D0 U9619 ( .A1(n24932), .A2(n3377), .B1(n25075), .B2(n4817), .C1(
        n24931), .C2(n3329), .ZN(n26753) );
  ND4D0 U9620 ( .A1(n26757), .A2(n26758), .A3(n26759), .A4(n26760), .ZN(n2175)
         );
  AN4D0 U9621 ( .A1(n26761), .A2(n26762), .A3(n26763), .A4(n26764), .Z(n26760)
         );
  NR4D0 U9622 ( .A1(n26765), .A2(n26766), .A3(n26767), .A4(n26768), .ZN(n26764) );
  OAI222D0 U9623 ( .A1(n24979), .A2(n15617), .B1(n24980), .B2(n4432), .C1(
        n24964), .C2(n2224), .ZN(n26768) );
  OAI222D0 U9624 ( .A1(n24920), .A2(n2512), .B1(n24981), .B2(n5152), .C1(
        n24963), .C2(n2416), .ZN(n26767) );
  OAI222D0 U9625 ( .A1(n24982), .A2(n4912), .B1(n24983), .B2(n4960), .C1(
        n24984), .C2(n4864), .ZN(n26766) );
  OAI222D0 U9626 ( .A1(n24985), .A2(n4384), .B1(n24986), .B2(n3760), .C1(
        n24987), .C2(n4336), .ZN(n26765) );
  NR4D0 U9627 ( .A1(n26769), .A2(n26770), .A3(n26771), .A4(n26772), .ZN(n26763) );
  OAI22D0 U9628 ( .A1(n24922), .A2(n2800), .B1(n24992), .B2(n3712), .ZN(n26772) );
  OAI222D0 U9629 ( .A1(n24993), .A2(n18052), .B1(n24962), .B2(n2752), .C1(
        n24994), .C2(n18053), .ZN(n26771) );
  OAI222D0 U9630 ( .A1(n24995), .A2(n5200), .B1(n24961), .B2(n2656), .C1(
        n24921), .C2(n2704), .ZN(n26770) );
  OAI222D0 U9631 ( .A1(n24927), .A2(n3136), .B1(n24996), .B2(n4768), .C1(
        n24997), .C2(n15616), .ZN(n26769) );
  NR4D0 U9632 ( .A1(n26773), .A2(n26774), .A3(n26775), .A4(n26776), .ZN(n26762) );
  OAI22D0 U9633 ( .A1(n24928), .A2(n3184), .B1(n24926), .B2(n3088), .ZN(n26776) );
  OAI222D0 U9634 ( .A1(n25002), .A2(n3424), .B1(n24929), .B2(n3232), .C1(
        n24933), .C2(n2320), .ZN(n26775) );
  OAI222D0 U9635 ( .A1(n25003), .A2(n3568), .B1(n25004), .B2(n3472), .C1(
        n25005), .C2(n3520), .ZN(n26774) );
  OAI222D0 U9636 ( .A1(n24965), .A2(n2560), .B1(n25006), .B2(n3616), .C1(
        n25007), .C2(n3664), .ZN(n26773) );
  NR4D0 U9637 ( .A1(n26777), .A2(n26778), .A3(n26779), .A4(n26780), .ZN(n26761) );
  OAI22D0 U9638 ( .A1(n25012), .A2(n5104), .B1(n24966), .B2(n2272), .ZN(n26780) );
  OAI222D0 U9639 ( .A1(n24925), .A2(n3040), .B1(n24923), .B2(n2944), .C1(
        n24960), .C2(n2848), .ZN(n26779) );
  OAI222D0 U9640 ( .A1(n25013), .A2(n5488), .B1(n25014), .B2(n5536), .C1(
        n24924), .C2(n2992), .ZN(n26778) );
  OAI222D0 U9641 ( .A1(n25015), .A2(n6064), .B1(n25016), .B2(n5968), .C1(
        n25017), .C2(n6112), .ZN(n26777) );
  INR4D0 U9642 ( .A1(n26781), .B1(n26782), .B2(n26783), .B3(n26784), .ZN(
        n26759) );
  OAI222D0 U9643 ( .A1(n25022), .A2(n5440), .B1(n25023), .B2(n6304), .C1(
        n25024), .C2(n5392), .ZN(n26784) );
  OAI222D0 U9644 ( .A1(n25025), .A2(n4480), .B1(n25026), .B2(n24685), .C1(
        n25027), .C2(n5584), .ZN(n26783) );
  OR4D0 U9645 ( .A1(n26785), .A2(n26786), .A3(n26787), .A4(n26788), .Z(n26782)
         );
  OAI222D0 U9646 ( .A1(n25032), .A2(n4576), .B1(n25033), .B2(n5296), .C1(
        n25034), .C2(n6208), .ZN(n26788) );
  OAI222D0 U9647 ( .A1(n25035), .A2(n6160), .B1(n25036), .B2(n4528), .C1(
        n25037), .C2(n5344), .ZN(n26787) );
  OAI22D0 U9648 ( .A1(n27207), .A2(n25038), .B1(n27206), .B2(n25039), .ZN(
        n26786) );
  OAI222D0 U9649 ( .A1(n24830), .A2(n25040), .B1(n25041), .B2(n5824), .C1(
        n25042), .C2(n5776), .ZN(n26785) );
  CKND0 U9650 ( .I(\Mem[44][42] ), .ZN(n24830) );
  AOI221D0 U9651 ( .A1(n27204), .A2(n25043), .B1(n27205), .B2(n25044), .C(
        n26789), .ZN(n26781) );
  OAI222D0 U9652 ( .A1(n25046), .A2(n6016), .B1(n24831), .B2(n25047), .C1(
        n25048), .C2(n4672), .ZN(n26789) );
  CKND0 U9653 ( .I(\Mem[45][42] ), .ZN(n24831) );
  NR4D0 U9654 ( .A1(n26790), .A2(n26791), .A3(n26792), .A4(n26793), .ZN(n26758) );
  OAI22D0 U9655 ( .A1(n25053), .A2(n5872), .B1(n25054), .B2(n5680), .ZN(n26793) );
  OAI222D0 U9656 ( .A1(n25055), .A2(n3808), .B1(n25056), .B2(n3856), .C1(
        n25057), .C2(n5920), .ZN(n26792) );
  OAI222D0 U9657 ( .A1(n25058), .A2(n3952), .B1(n25059), .B2(n4000), .C1(
        n25060), .C2(n3904), .ZN(n26791) );
  OAI222D0 U9658 ( .A1(n25061), .A2(n4096), .B1(n25062), .B2(n4144), .C1(
        n25063), .C2(n4048), .ZN(n26790) );
  NR4D0 U9659 ( .A1(n26794), .A2(n26795), .A3(n26796), .A4(n26797), .ZN(n26757) );
  OAI22D0 U9660 ( .A1(n25068), .A2(n2368), .B1(n25069), .B2(n2896), .ZN(n26797) );
  OAI222D0 U9661 ( .A1(n25070), .A2(n2464), .B1(n25071), .B2(n4288), .C1(
        n25072), .C2(n2608), .ZN(n26796) );
  OAI222D0 U9662 ( .A1(n25073), .A2(n4240), .B1(n24930), .B2(n3280), .C1(
        n25074), .C2(n4192), .ZN(n26795) );
  OAI222D0 U9663 ( .A1(n24932), .A2(n3376), .B1(n25075), .B2(n4816), .C1(
        n24931), .C2(n3328), .ZN(n26794) );
  ND4D0 U9664 ( .A1(n26798), .A2(n26799), .A3(n26800), .A4(n26801), .ZN(n2174)
         );
  AN4D0 U9665 ( .A1(n26802), .A2(n26803), .A3(n26804), .A4(n26805), .Z(n26801)
         );
  NR4D0 U9666 ( .A1(n26806), .A2(n26807), .A3(n26808), .A4(n26809), .ZN(n26805) );
  OAI222D0 U9667 ( .A1(n24979), .A2(n15621), .B1(n24980), .B2(n4431), .C1(
        n24964), .C2(n2223), .ZN(n26809) );
  OAI222D0 U9668 ( .A1(n24920), .A2(n2511), .B1(n24981), .B2(n5151), .C1(
        n24963), .C2(n2415), .ZN(n26808) );
  OAI222D0 U9669 ( .A1(n24982), .A2(n4911), .B1(n24983), .B2(n4959), .C1(
        n24984), .C2(n4863), .ZN(n26807) );
  OAI222D0 U9670 ( .A1(n24985), .A2(n4383), .B1(n24986), .B2(n3759), .C1(
        n24987), .C2(n4335), .ZN(n26806) );
  NR4D0 U9671 ( .A1(n26810), .A2(n26811), .A3(n26812), .A4(n26813), .ZN(n26804) );
  OAI22D0 U9672 ( .A1(n24922), .A2(n2799), .B1(n24992), .B2(n3711), .ZN(n26813) );
  OAI222D0 U9673 ( .A1(n24993), .A2(n18055), .B1(n24962), .B2(n2751), .C1(
        n24994), .C2(n18056), .ZN(n26812) );
  OAI222D0 U9674 ( .A1(n24995), .A2(n5199), .B1(n24961), .B2(n2655), .C1(
        n24921), .C2(n2703), .ZN(n26811) );
  OAI222D0 U9675 ( .A1(n24927), .A2(n3135), .B1(n24996), .B2(n4767), .C1(
        n24997), .C2(n15620), .ZN(n26810) );
  NR4D0 U9676 ( .A1(n26814), .A2(n26815), .A3(n26816), .A4(n26817), .ZN(n26803) );
  OAI22D0 U9677 ( .A1(n24928), .A2(n3183), .B1(n24926), .B2(n3087), .ZN(n26817) );
  OAI222D0 U9678 ( .A1(n25002), .A2(n3423), .B1(n24929), .B2(n3231), .C1(
        n24933), .C2(n2319), .ZN(n26816) );
  OAI222D0 U9679 ( .A1(n25003), .A2(n3567), .B1(n25004), .B2(n3471), .C1(
        n25005), .C2(n3519), .ZN(n26815) );
  OAI222D0 U9680 ( .A1(n24965), .A2(n2559), .B1(n25006), .B2(n3615), .C1(
        n25007), .C2(n3663), .ZN(n26814) );
  NR4D0 U9681 ( .A1(n26818), .A2(n26819), .A3(n26820), .A4(n26821), .ZN(n26802) );
  OAI22D0 U9682 ( .A1(n25012), .A2(n5103), .B1(n24966), .B2(n2271), .ZN(n26821) );
  OAI222D0 U9683 ( .A1(n24925), .A2(n3039), .B1(n24923), .B2(n2943), .C1(
        n24960), .C2(n2847), .ZN(n26820) );
  OAI222D0 U9684 ( .A1(n25013), .A2(n5487), .B1(n25014), .B2(n5535), .C1(
        n24924), .C2(n2991), .ZN(n26819) );
  OAI222D0 U9685 ( .A1(n25015), .A2(n6063), .B1(n25016), .B2(n5967), .C1(
        n25017), .C2(n6111), .ZN(n26818) );
  INR4D0 U9686 ( .A1(n26822), .B1(n26823), .B2(n26824), .B3(n26825), .ZN(
        n26800) );
  OAI222D0 U9687 ( .A1(n25022), .A2(n5439), .B1(n25023), .B2(n6303), .C1(
        n25024), .C2(n5391), .ZN(n26825) );
  OAI222D0 U9688 ( .A1(n25025), .A2(n4479), .B1(n25026), .B2(n24688), .C1(
        n25027), .C2(n5583), .ZN(n26824) );
  OR4D0 U9689 ( .A1(n26826), .A2(n26827), .A3(n26828), .A4(n26829), .Z(n26823)
         );
  OAI222D0 U9690 ( .A1(n25032), .A2(n4575), .B1(n25033), .B2(n5295), .C1(
        n25034), .C2(n6207), .ZN(n26829) );
  OAI222D0 U9691 ( .A1(n25035), .A2(n6159), .B1(n25036), .B2(n4527), .C1(
        n25037), .C2(n5343), .ZN(n26828) );
  OAI22D0 U9692 ( .A1(n27211), .A2(n25038), .B1(n27210), .B2(n25039), .ZN(
        n26827) );
  OAI222D0 U9693 ( .A1(n24828), .A2(n25040), .B1(n25041), .B2(n5823), .C1(
        n25042), .C2(n5775), .ZN(n26826) );
  CKND0 U9694 ( .I(\Mem[44][43] ), .ZN(n24828) );
  AOI221D0 U9695 ( .A1(n27208), .A2(n25043), .B1(n27209), .B2(n25044), .C(
        n26830), .ZN(n26822) );
  OAI222D0 U9696 ( .A1(n25046), .A2(n6015), .B1(n24829), .B2(n25047), .C1(
        n25048), .C2(n4671), .ZN(n26830) );
  CKND0 U9697 ( .I(\Mem[45][43] ), .ZN(n24829) );
  NR4D0 U9698 ( .A1(n26831), .A2(n26832), .A3(n26833), .A4(n26834), .ZN(n26799) );
  OAI22D0 U9699 ( .A1(n25053), .A2(n5871), .B1(n25054), .B2(n5679), .ZN(n26834) );
  OAI222D0 U9700 ( .A1(n25055), .A2(n3807), .B1(n25056), .B2(n3855), .C1(
        n25057), .C2(n5919), .ZN(n26833) );
  OAI222D0 U9701 ( .A1(n25058), .A2(n3951), .B1(n25059), .B2(n3999), .C1(
        n25060), .C2(n3903), .ZN(n26832) );
  OAI222D0 U9702 ( .A1(n25061), .A2(n4095), .B1(n25062), .B2(n4143), .C1(
        n25063), .C2(n4047), .ZN(n26831) );
  NR4D0 U9703 ( .A1(n26835), .A2(n26836), .A3(n26837), .A4(n26838), .ZN(n26798) );
  OAI22D0 U9704 ( .A1(n25068), .A2(n2367), .B1(n25069), .B2(n2895), .ZN(n26838) );
  OAI222D0 U9705 ( .A1(n25070), .A2(n2463), .B1(n25071), .B2(n4287), .C1(
        n25072), .C2(n2607), .ZN(n26837) );
  OAI222D0 U9706 ( .A1(n25073), .A2(n4239), .B1(n24930), .B2(n3279), .C1(
        n25074), .C2(n4191), .ZN(n26836) );
  OAI222D0 U9707 ( .A1(n24932), .A2(n3375), .B1(n25075), .B2(n4815), .C1(
        n24931), .C2(n3327), .ZN(n26835) );
  ND4D0 U9708 ( .A1(n26839), .A2(n26840), .A3(n26841), .A4(n26842), .ZN(n2173)
         );
  AN4D0 U9709 ( .A1(n26843), .A2(n26844), .A3(n26845), .A4(n26846), .Z(n26842)
         );
  NR4D0 U9710 ( .A1(n26847), .A2(n26848), .A3(n26849), .A4(n26850), .ZN(n26846) );
  OAI222D0 U9711 ( .A1(n24979), .A2(n15625), .B1(n24980), .B2(n4430), .C1(
        n24964), .C2(n2222), .ZN(n26850) );
  OAI222D0 U9712 ( .A1(n24920), .A2(n2510), .B1(n24981), .B2(n5150), .C1(
        n24963), .C2(n2414), .ZN(n26849) );
  OAI222D0 U9713 ( .A1(n24982), .A2(n4910), .B1(n24983), .B2(n4958), .C1(
        n24984), .C2(n4862), .ZN(n26848) );
  OAI222D0 U9714 ( .A1(n24985), .A2(n4382), .B1(n24986), .B2(n3758), .C1(
        n24987), .C2(n4334), .ZN(n26847) );
  NR4D0 U9715 ( .A1(n26851), .A2(n26852), .A3(n26853), .A4(n26854), .ZN(n26845) );
  OAI22D0 U9716 ( .A1(n24922), .A2(n2798), .B1(n24992), .B2(n3710), .ZN(n26854) );
  OAI222D0 U9717 ( .A1(n24993), .A2(n18058), .B1(n24962), .B2(n2750), .C1(
        n24994), .C2(n18059), .ZN(n26853) );
  OAI222D0 U9718 ( .A1(n24995), .A2(n5198), .B1(n24961), .B2(n2654), .C1(
        n24921), .C2(n2702), .ZN(n26852) );
  OAI222D0 U9719 ( .A1(n24927), .A2(n3134), .B1(n24996), .B2(n4766), .C1(
        n24997), .C2(n15624), .ZN(n26851) );
  NR4D0 U9720 ( .A1(n26855), .A2(n26856), .A3(n26857), .A4(n26858), .ZN(n26844) );
  OAI22D0 U9721 ( .A1(n24928), .A2(n3182), .B1(n24926), .B2(n3086), .ZN(n26858) );
  OAI222D0 U9722 ( .A1(n25002), .A2(n3422), .B1(n24929), .B2(n3230), .C1(
        n24933), .C2(n2318), .ZN(n26857) );
  OAI222D0 U9723 ( .A1(n25003), .A2(n3566), .B1(n25004), .B2(n3470), .C1(
        n25005), .C2(n3518), .ZN(n26856) );
  OAI222D0 U9724 ( .A1(n24965), .A2(n2558), .B1(n25006), .B2(n3614), .C1(
        n25007), .C2(n3662), .ZN(n26855) );
  NR4D0 U9725 ( .A1(n26859), .A2(n26860), .A3(n26861), .A4(n26862), .ZN(n26843) );
  OAI22D0 U9726 ( .A1(n25012), .A2(n5102), .B1(n24966), .B2(n2270), .ZN(n26862) );
  OAI222D0 U9727 ( .A1(n24925), .A2(n3038), .B1(n24923), .B2(n2942), .C1(
        n24960), .C2(n2846), .ZN(n26861) );
  OAI222D0 U9728 ( .A1(n25013), .A2(n5486), .B1(n25014), .B2(n5534), .C1(
        n24924), .C2(n2990), .ZN(n26860) );
  OAI222D0 U9729 ( .A1(n25015), .A2(n6062), .B1(n25016), .B2(n5966), .C1(
        n25017), .C2(n6110), .ZN(n26859) );
  INR4D0 U9730 ( .A1(n26863), .B1(n26864), .B2(n26865), .B3(n26866), .ZN(
        n26841) );
  OAI222D0 U9731 ( .A1(n25022), .A2(n5438), .B1(n25023), .B2(n6302), .C1(
        n25024), .C2(n5390), .ZN(n26866) );
  OAI222D0 U9732 ( .A1(n25025), .A2(n4478), .B1(n25026), .B2(n24691), .C1(
        n25027), .C2(n5582), .ZN(n26865) );
  OR4D0 U9733 ( .A1(n26867), .A2(n26868), .A3(n26869), .A4(n26870), .Z(n26864)
         );
  OAI222D0 U9734 ( .A1(n25032), .A2(n4574), .B1(n25033), .B2(n5294), .C1(
        n25034), .C2(n6206), .ZN(n26870) );
  OAI222D0 U9735 ( .A1(n25035), .A2(n6158), .B1(n25036), .B2(n4526), .C1(
        n25037), .C2(n5342), .ZN(n26869) );
  OAI22D0 U9736 ( .A1(n27215), .A2(n25038), .B1(n27214), .B2(n25039), .ZN(
        n26868) );
  OAI222D0 U9737 ( .A1(n24826), .A2(n25040), .B1(n25041), .B2(n5822), .C1(
        n25042), .C2(n5774), .ZN(n26867) );
  CKND0 U9738 ( .I(\Mem[44][44] ), .ZN(n24826) );
  AOI221D0 U9739 ( .A1(n27212), .A2(n25043), .B1(n27213), .B2(n25044), .C(
        n26871), .ZN(n26863) );
  OAI222D0 U9740 ( .A1(n25046), .A2(n6014), .B1(n24827), .B2(n25047), .C1(
        n25048), .C2(n4670), .ZN(n26871) );
  CKND0 U9741 ( .I(\Mem[45][44] ), .ZN(n24827) );
  NR4D0 U9742 ( .A1(n26872), .A2(n26873), .A3(n26874), .A4(n26875), .ZN(n26840) );
  OAI22D0 U9743 ( .A1(n25053), .A2(n5870), .B1(n25054), .B2(n5678), .ZN(n26875) );
  OAI222D0 U9744 ( .A1(n25055), .A2(n3806), .B1(n25056), .B2(n3854), .C1(
        n25057), .C2(n5918), .ZN(n26874) );
  OAI222D0 U9745 ( .A1(n25058), .A2(n3950), .B1(n25059), .B2(n3998), .C1(
        n25060), .C2(n3902), .ZN(n26873) );
  OAI222D0 U9746 ( .A1(n25061), .A2(n4094), .B1(n25062), .B2(n4142), .C1(
        n25063), .C2(n4046), .ZN(n26872) );
  NR4D0 U9747 ( .A1(n26876), .A2(n26877), .A3(n26878), .A4(n26879), .ZN(n26839) );
  OAI22D0 U9748 ( .A1(n25068), .A2(n2366), .B1(n25069), .B2(n2894), .ZN(n26879) );
  OAI222D0 U9749 ( .A1(n25070), .A2(n2462), .B1(n25071), .B2(n4286), .C1(
        n25072), .C2(n2606), .ZN(n26878) );
  OAI222D0 U9750 ( .A1(n25073), .A2(n4238), .B1(n24930), .B2(n3278), .C1(
        n25074), .C2(n4190), .ZN(n26877) );
  OAI222D0 U9751 ( .A1(n24932), .A2(n3374), .B1(n25075), .B2(n4814), .C1(
        n24931), .C2(n3326), .ZN(n26876) );
  ND4D0 U9752 ( .A1(n26880), .A2(n26881), .A3(n26882), .A4(n26883), .ZN(n2172)
         );
  AN4D0 U9753 ( .A1(n26884), .A2(n26885), .A3(n26886), .A4(n26887), .Z(n26883)
         );
  NR4D0 U9754 ( .A1(n26888), .A2(n26889), .A3(n26890), .A4(n26891), .ZN(n26887) );
  OAI222D0 U9755 ( .A1(n24979), .A2(n15629), .B1(n24980), .B2(n4429), .C1(
        n24964), .C2(n2221), .ZN(n26891) );
  OAI222D0 U9756 ( .A1(n24920), .A2(n2509), .B1(n24981), .B2(n5149), .C1(
        n24963), .C2(n2413), .ZN(n26890) );
  OAI222D0 U9757 ( .A1(n24982), .A2(n4909), .B1(n24983), .B2(n4957), .C1(
        n24984), .C2(n4861), .ZN(n26889) );
  OAI222D0 U9758 ( .A1(n24985), .A2(n4381), .B1(n24986), .B2(n3757), .C1(
        n24987), .C2(n4333), .ZN(n26888) );
  NR4D0 U9759 ( .A1(n26892), .A2(n26893), .A3(n26894), .A4(n26895), .ZN(n26886) );
  OAI22D0 U9760 ( .A1(n24922), .A2(n2797), .B1(n24992), .B2(n3709), .ZN(n26895) );
  OAI222D0 U9761 ( .A1(n24993), .A2(n18061), .B1(n24962), .B2(n2749), .C1(
        n24994), .C2(n18062), .ZN(n26894) );
  OAI222D0 U9762 ( .A1(n24995), .A2(n5197), .B1(n24961), .B2(n2653), .C1(
        n24921), .C2(n2701), .ZN(n26893) );
  OAI222D0 U9763 ( .A1(n24927), .A2(n3133), .B1(n24996), .B2(n4765), .C1(
        n24997), .C2(n15628), .ZN(n26892) );
  NR4D0 U9764 ( .A1(n26896), .A2(n26897), .A3(n26898), .A4(n26899), .ZN(n26885) );
  OAI22D0 U9765 ( .A1(n24928), .A2(n3181), .B1(n24926), .B2(n3085), .ZN(n26899) );
  OAI222D0 U9766 ( .A1(n25002), .A2(n3421), .B1(n24929), .B2(n3229), .C1(
        n24933), .C2(n2317), .ZN(n26898) );
  OAI222D0 U9767 ( .A1(n25003), .A2(n3565), .B1(n25004), .B2(n3469), .C1(
        n25005), .C2(n3517), .ZN(n26897) );
  OAI222D0 U9768 ( .A1(n24965), .A2(n2557), .B1(n25006), .B2(n3613), .C1(
        n25007), .C2(n3661), .ZN(n26896) );
  NR4D0 U9769 ( .A1(n26900), .A2(n26901), .A3(n26902), .A4(n26903), .ZN(n26884) );
  OAI22D0 U9770 ( .A1(n25012), .A2(n5101), .B1(n24966), .B2(n2269), .ZN(n26903) );
  OAI222D0 U9771 ( .A1(n24925), .A2(n3037), .B1(n24923), .B2(n2941), .C1(
        n24960), .C2(n2845), .ZN(n26902) );
  OAI222D0 U9772 ( .A1(n25013), .A2(n5485), .B1(n25014), .B2(n5533), .C1(
        n24924), .C2(n2989), .ZN(n26901) );
  OAI222D0 U9773 ( .A1(n25015), .A2(n6061), .B1(n25016), .B2(n5965), .C1(
        n25017), .C2(n6109), .ZN(n26900) );
  INR4D0 U9774 ( .A1(n26904), .B1(n26905), .B2(n26906), .B3(n26907), .ZN(
        n26882) );
  OAI222D0 U9775 ( .A1(n25022), .A2(n5437), .B1(n25023), .B2(n6301), .C1(
        n25024), .C2(n5389), .ZN(n26907) );
  OAI222D0 U9776 ( .A1(n25025), .A2(n4477), .B1(n25026), .B2(n24694), .C1(
        n25027), .C2(n5581), .ZN(n26906) );
  OR4D0 U9777 ( .A1(n26908), .A2(n26909), .A3(n26910), .A4(n26911), .Z(n26905)
         );
  OAI222D0 U9778 ( .A1(n25032), .A2(n4573), .B1(n25033), .B2(n5293), .C1(
        n25034), .C2(n6205), .ZN(n26911) );
  OAI222D0 U9779 ( .A1(n25035), .A2(n6157), .B1(n25036), .B2(n4525), .C1(
        n25037), .C2(n5341), .ZN(n26910) );
  OAI22D0 U9780 ( .A1(n27219), .A2(n25038), .B1(n27218), .B2(n25039), .ZN(
        n26909) );
  OAI222D0 U9781 ( .A1(n24824), .A2(n25040), .B1(n25041), .B2(n5821), .C1(
        n25042), .C2(n5773), .ZN(n26908) );
  CKND0 U9782 ( .I(\Mem[44][45] ), .ZN(n24824) );
  AOI221D0 U9783 ( .A1(n27216), .A2(n25043), .B1(n27217), .B2(n25044), .C(
        n26912), .ZN(n26904) );
  OAI222D0 U9784 ( .A1(n25046), .A2(n6013), .B1(n24825), .B2(n25047), .C1(
        n25048), .C2(n4669), .ZN(n26912) );
  CKND0 U9785 ( .I(\Mem[45][45] ), .ZN(n24825) );
  NR4D0 U9786 ( .A1(n26913), .A2(n26914), .A3(n26915), .A4(n26916), .ZN(n26881) );
  OAI22D0 U9787 ( .A1(n25053), .A2(n5869), .B1(n25054), .B2(n5677), .ZN(n26916) );
  OAI222D0 U9788 ( .A1(n25055), .A2(n3805), .B1(n25056), .B2(n3853), .C1(
        n25057), .C2(n5917), .ZN(n26915) );
  OAI222D0 U9789 ( .A1(n25058), .A2(n3949), .B1(n25059), .B2(n3997), .C1(
        n25060), .C2(n3901), .ZN(n26914) );
  OAI222D0 U9790 ( .A1(n25061), .A2(n4093), .B1(n25062), .B2(n4141), .C1(
        n25063), .C2(n4045), .ZN(n26913) );
  NR4D0 U9791 ( .A1(n26917), .A2(n26918), .A3(n26919), .A4(n26920), .ZN(n26880) );
  OAI22D0 U9792 ( .A1(n25068), .A2(n2365), .B1(n25069), .B2(n2893), .ZN(n26920) );
  OAI222D0 U9793 ( .A1(n25070), .A2(n2461), .B1(n25071), .B2(n4285), .C1(
        n25072), .C2(n2605), .ZN(n26919) );
  OAI222D0 U9794 ( .A1(n25073), .A2(n4237), .B1(n24930), .B2(n3277), .C1(
        n25074), .C2(n4189), .ZN(n26918) );
  OAI222D0 U9795 ( .A1(n24932), .A2(n3373), .B1(n25075), .B2(n4813), .C1(
        n24931), .C2(n3325), .ZN(n26917) );
  ND4D0 U9796 ( .A1(n26921), .A2(n26922), .A3(n26923), .A4(n26924), .ZN(n2171)
         );
  AN4D0 U9797 ( .A1(n26925), .A2(n26926), .A3(n26927), .A4(n26928), .Z(n26924)
         );
  NR4D0 U9798 ( .A1(n26929), .A2(n26930), .A3(n26931), .A4(n26932), .ZN(n26928) );
  OAI222D0 U9799 ( .A1(n24979), .A2(n15633), .B1(n24980), .B2(n4428), .C1(
        n24964), .C2(n2220), .ZN(n26932) );
  OAI222D0 U9800 ( .A1(n24920), .A2(n2508), .B1(n24981), .B2(n5148), .C1(
        n24963), .C2(n2412), .ZN(n26931) );
  OAI222D0 U9801 ( .A1(n24982), .A2(n4908), .B1(n24983), .B2(n4956), .C1(
        n24984), .C2(n4860), .ZN(n26930) );
  OAI222D0 U9802 ( .A1(n24985), .A2(n4380), .B1(n24986), .B2(n3756), .C1(
        n24987), .C2(n4332), .ZN(n26929) );
  NR4D0 U9803 ( .A1(n26933), .A2(n26934), .A3(n26935), .A4(n26936), .ZN(n26927) );
  OAI22D0 U9804 ( .A1(n24922), .A2(n2796), .B1(n24992), .B2(n3708), .ZN(n26936) );
  OAI222D0 U9805 ( .A1(n24993), .A2(n18064), .B1(n24962), .B2(n2748), .C1(
        n24994), .C2(n18065), .ZN(n26935) );
  OAI222D0 U9806 ( .A1(n24995), .A2(n5196), .B1(n24961), .B2(n2652), .C1(
        n24921), .C2(n2700), .ZN(n26934) );
  OAI222D0 U9807 ( .A1(n24927), .A2(n3132), .B1(n24996), .B2(n4764), .C1(
        n24997), .C2(n15632), .ZN(n26933) );
  NR4D0 U9808 ( .A1(n26937), .A2(n26938), .A3(n26939), .A4(n26940), .ZN(n26926) );
  OAI22D0 U9809 ( .A1(n24928), .A2(n3180), .B1(n24926), .B2(n3084), .ZN(n26940) );
  OAI222D0 U9810 ( .A1(n25002), .A2(n3420), .B1(n24929), .B2(n3228), .C1(
        n24933), .C2(n2316), .ZN(n26939) );
  OAI222D0 U9811 ( .A1(n25003), .A2(n3564), .B1(n25004), .B2(n3468), .C1(
        n25005), .C2(n3516), .ZN(n26938) );
  OAI222D0 U9812 ( .A1(n24965), .A2(n2556), .B1(n25006), .B2(n3612), .C1(
        n25007), .C2(n3660), .ZN(n26937) );
  NR4D0 U9813 ( .A1(n26941), .A2(n26942), .A3(n26943), .A4(n26944), .ZN(n26925) );
  OAI22D0 U9814 ( .A1(n25012), .A2(n5100), .B1(n24966), .B2(n2268), .ZN(n26944) );
  OAI222D0 U9815 ( .A1(n24925), .A2(n3036), .B1(n24923), .B2(n2940), .C1(
        n24960), .C2(n2844), .ZN(n26943) );
  OAI222D0 U9816 ( .A1(n25013), .A2(n5484), .B1(n25014), .B2(n5532), .C1(
        n24924), .C2(n2988), .ZN(n26942) );
  OAI222D0 U9817 ( .A1(n25015), .A2(n6060), .B1(n25016), .B2(n5964), .C1(
        n25017), .C2(n6108), .ZN(n26941) );
  INR4D0 U9818 ( .A1(n26945), .B1(n26946), .B2(n26947), .B3(n26948), .ZN(
        n26923) );
  OAI222D0 U9819 ( .A1(n25022), .A2(n5436), .B1(n25023), .B2(n6300), .C1(
        n25024), .C2(n5388), .ZN(n26948) );
  OAI222D0 U9820 ( .A1(n25025), .A2(n4476), .B1(n25026), .B2(n24697), .C1(
        n25027), .C2(n5580), .ZN(n26947) );
  OR4D0 U9821 ( .A1(n26949), .A2(n26950), .A3(n26951), .A4(n26952), .Z(n26946)
         );
  OAI222D0 U9822 ( .A1(n25032), .A2(n4572), .B1(n25033), .B2(n5292), .C1(
        n25034), .C2(n6204), .ZN(n26952) );
  OAI222D0 U9823 ( .A1(n25035), .A2(n6156), .B1(n25036), .B2(n4524), .C1(
        n25037), .C2(n5340), .ZN(n26951) );
  OAI22D0 U9824 ( .A1(n27223), .A2(n25038), .B1(n27222), .B2(n25039), .ZN(
        n26950) );
  OAI222D0 U9825 ( .A1(n24822), .A2(n25040), .B1(n25041), .B2(n5820), .C1(
        n25042), .C2(n5772), .ZN(n26949) );
  CKND0 U9826 ( .I(\Mem[44][46] ), .ZN(n24822) );
  AOI221D0 U9827 ( .A1(n27220), .A2(n25043), .B1(n27221), .B2(n25044), .C(
        n26953), .ZN(n26945) );
  OAI222D0 U9828 ( .A1(n25046), .A2(n6012), .B1(n24823), .B2(n25047), .C1(
        n25048), .C2(n4668), .ZN(n26953) );
  CKND0 U9829 ( .I(\Mem[45][46] ), .ZN(n24823) );
  NR4D0 U9830 ( .A1(n26954), .A2(n26955), .A3(n26956), .A4(n26957), .ZN(n26922) );
  OAI22D0 U9831 ( .A1(n25053), .A2(n5868), .B1(n25054), .B2(n5676), .ZN(n26957) );
  OAI222D0 U9832 ( .A1(n25055), .A2(n3804), .B1(n25056), .B2(n3852), .C1(
        n25057), .C2(n5916), .ZN(n26956) );
  OAI222D0 U9833 ( .A1(n25058), .A2(n3948), .B1(n25059), .B2(n3996), .C1(
        n25060), .C2(n3900), .ZN(n26955) );
  OAI222D0 U9834 ( .A1(n25061), .A2(n4092), .B1(n25062), .B2(n4140), .C1(
        n25063), .C2(n4044), .ZN(n26954) );
  NR4D0 U9835 ( .A1(n26958), .A2(n26959), .A3(n26960), .A4(n26961), .ZN(n26921) );
  OAI22D0 U9836 ( .A1(n25068), .A2(n2364), .B1(n25069), .B2(n2892), .ZN(n26961) );
  OAI222D0 U9837 ( .A1(n25070), .A2(n2460), .B1(n25071), .B2(n4284), .C1(
        n25072), .C2(n2604), .ZN(n26960) );
  OAI222D0 U9838 ( .A1(n25073), .A2(n4236), .B1(n24930), .B2(n3276), .C1(
        n25074), .C2(n4188), .ZN(n26959) );
  OAI222D0 U9839 ( .A1(n24932), .A2(n3372), .B1(n25075), .B2(n4812), .C1(
        n24931), .C2(n3324), .ZN(n26958) );
  ND4D0 U9840 ( .A1(n26962), .A2(n26963), .A3(n26964), .A4(n26965), .ZN(n2170)
         );
  AN4D0 U9841 ( .A1(n26966), .A2(n26967), .A3(n26968), .A4(n26969), .Z(n26965)
         );
  NR4D0 U9842 ( .A1(n26970), .A2(n26971), .A3(n26972), .A4(n26973), .ZN(n26969) );
  OAI222D0 U9843 ( .A1(n24979), .A2(n15637), .B1(n24980), .B2(n4427), .C1(
        n24964), .C2(n2219), .ZN(n26973) );
  CKND2D0 U9844 ( .A1(n24959), .A2(n26976), .ZN(n24979) );
  OAI222D0 U9845 ( .A1(n24920), .A2(n2507), .B1(n24981), .B2(n5147), .C1(
        n24963), .C2(n2411), .ZN(n26972) );
  OAI222D0 U9846 ( .A1(n24982), .A2(n4907), .B1(n24983), .B2(n4955), .C1(
        n24984), .C2(n4859), .ZN(n26971) );
  CKND2D0 U9847 ( .A1(n24951), .A2(n26982), .ZN(n24982) );
  OAI222D0 U9848 ( .A1(n24985), .A2(n4379), .B1(n24986), .B2(n3755), .C1(
        n24987), .C2(n4331), .ZN(n26970) );
  CKND2D0 U9849 ( .A1(n26978), .A2(n24952), .ZN(n24985) );
  NR4D0 U9850 ( .A1(n26984), .A2(n26985), .A3(n26986), .A4(n26987), .ZN(n26968) );
  OAI22D0 U9851 ( .A1(n24922), .A2(n2795), .B1(n24992), .B2(n3707), .ZN(n26987) );
  CKND2D0 U9852 ( .A1(n26988), .A2(n26978), .ZN(n24992) );
  OAI222D0 U9853 ( .A1(n24993), .A2(n18067), .B1(n24962), .B2(n2747), .C1(
        n24994), .C2(n18068), .ZN(n26986) );
  CKND2D0 U9854 ( .A1(n24951), .A2(n26989), .ZN(n24993) );
  OAI222D0 U9855 ( .A1(n24995), .A2(n5195), .B1(n24961), .B2(n2651), .C1(
        n24921), .C2(n2699), .ZN(n26985) );
  CKND2D0 U9856 ( .A1(n24959), .A2(n26974), .ZN(n24995) );
  OAI222D0 U9857 ( .A1(n24927), .A2(n3131), .B1(n24996), .B2(n4763), .C1(
        n24997), .C2(n15636), .ZN(n26984) );
  NR4D0 U9858 ( .A1(n26993), .A2(n26994), .A3(n26995), .A4(n26996), .ZN(n26967) );
  OAI22D0 U9859 ( .A1(n24928), .A2(n3179), .B1(n24926), .B2(n3083), .ZN(n26996) );
  OAI222D0 U9860 ( .A1(n25002), .A2(n3419), .B1(n24929), .B2(n3227), .C1(
        n24933), .C2(n2315), .ZN(n26995) );
  CKND2D0 U9861 ( .A1(n26980), .A2(n26988), .ZN(n25002) );
  OAI222D0 U9862 ( .A1(n25003), .A2(n3563), .B1(n25004), .B2(n3467), .C1(
        n25005), .C2(n3515), .ZN(n26994) );
  CKND2D0 U9863 ( .A1(n26988), .A2(n26989), .ZN(n25003) );
  OAI222D0 U9864 ( .A1(n24965), .A2(n2555), .B1(n25006), .B2(n3611), .C1(
        n25007), .C2(n3659), .ZN(n26993) );
  NR4D0 U9865 ( .A1(n26999), .A2(n27000), .A3(n27001), .A4(n27002), .ZN(n26966) );
  OAI22D0 U9866 ( .A1(n25012), .A2(n5099), .B1(n24966), .B2(n2267), .ZN(n27002) );
  CKND2D0 U9867 ( .A1(n26983), .A2(n24951), .ZN(n25012) );
  OAI222D0 U9868 ( .A1(n24925), .A2(n3035), .B1(n24923), .B2(n2939), .C1(
        n24960), .C2(n2843), .ZN(n27001) );
  OAI222D0 U9869 ( .A1(n25013), .A2(n5483), .B1(n25014), .B2(n5531), .C1(
        n24924), .C2(n2987), .ZN(n27000) );
  CKND2D0 U9870 ( .A1(n24959), .A2(n26979), .ZN(n25013) );
  OAI222D0 U9871 ( .A1(n25015), .A2(n6059), .B1(n25016), .B2(n5963), .C1(
        n25017), .C2(n6107), .ZN(n26999) );
  CKND0 U9872 ( .I(n24948), .ZN(n26974) );
  CKND2D0 U9873 ( .A1(n27005), .A2(n27006), .ZN(n24948) );
  CKND2D0 U9874 ( .A1(n27007), .A2(n27004), .ZN(n25015) );
  INR4D0 U9875 ( .A1(n27008), .B1(n27009), .B2(n27010), .B3(n27011), .ZN(
        n26964) );
  OAI222D0 U9876 ( .A1(n25022), .A2(n5435), .B1(n25023), .B2(n6299), .C1(
        n25024), .C2(n5387), .ZN(n27011) );
  CKND2D0 U9877 ( .A1(n24959), .A2(n26998), .ZN(n25022) );
  OAI222D0 U9878 ( .A1(n25025), .A2(n4475), .B1(n25026), .B2(n24700), .C1(
        n25027), .C2(n5579), .ZN(n27010) );
  CKND2D0 U9879 ( .A1(n24951), .A2(n26976), .ZN(n25025) );
  OR4D0 U9880 ( .A1(n27014), .A2(n27015), .A3(n27016), .A4(n27017), .Z(n27009)
         );
  OAI222D0 U9881 ( .A1(n25032), .A2(n4571), .B1(n25033), .B2(n5291), .C1(
        n25034), .C2(n6203), .ZN(n27017) );
  CKND2D0 U9882 ( .A1(n24951), .A2(n26992), .ZN(n25032) );
  OAI222D0 U9883 ( .A1(n25035), .A2(n6155), .B1(n25036), .B2(n4523), .C1(
        n25037), .C2(n5339), .ZN(n27016) );
  NR2D0 U9884 ( .A1(n24950), .A2(Address[4]), .ZN(n24959) );
  CKND2D0 U9885 ( .A1(n27007), .A2(n27018), .ZN(n25035) );
  AN2D0 U9886 ( .A1(n24957), .A2(n27019), .Z(n27007) );
  OAI22D0 U9887 ( .A1(n27227), .A2(n25038), .B1(n27226), .B2(n25039), .ZN(
        n27015) );
  OAI222D0 U9888 ( .A1(n24818), .A2(n25040), .B1(n25041), .B2(n5819), .C1(
        n25042), .C2(n5771), .ZN(n27014) );
  CKND2D0 U9889 ( .A1(n27018), .A2(n27020), .ZN(n24915) );
  CKND0 U9890 ( .I(\Mem[44][47] ), .ZN(n24818) );
  AOI221D0 U9891 ( .A1(n27224), .A2(n25043), .B1(n27225), .B2(n25044), .C(
        n27021), .ZN(n27008) );
  OAI222D0 U9892 ( .A1(n25046), .A2(n6011), .B1(n24820), .B2(n25047), .C1(
        n25048), .C2(n4667), .ZN(n27021) );
  CKND0 U9893 ( .I(n24918), .ZN(n26990) );
  CKND2D0 U9894 ( .A1(n27022), .A2(n27018), .ZN(n24918) );
  CKND0 U9895 ( .I(\Mem[45][47] ), .ZN(n24820) );
  CKND2D0 U9896 ( .A1(n27003), .A2(n27005), .ZN(n25046) );
  AN2D0 U9897 ( .A1(n24957), .A2(Address[0]), .Z(n27003) );
  AN2D0 U9898 ( .A1(n24951), .A2(n26977), .Z(n25043) );
  NR4D0 U9899 ( .A1(n27024), .A2(n27025), .A3(n27026), .A4(n27027), .ZN(n26963) );
  OAI22D0 U9900 ( .A1(n25053), .A2(n5867), .B1(n25054), .B2(n5675), .ZN(n27027) );
  CKND2D0 U9901 ( .A1(Address[6]), .A2(n26982), .ZN(n25054) );
  CKND2D0 U9902 ( .A1(Address[6]), .A2(n26983), .ZN(n25053) );
  OAI222D0 U9903 ( .A1(n25055), .A2(n3803), .B1(n25056), .B2(n3851), .C1(
        n25057), .C2(n5915), .ZN(n27026) );
  CKND2D0 U9904 ( .A1(n27012), .A2(n27022), .ZN(n24934) );
  CKND2D0 U9905 ( .A1(n27004), .A2(n27006), .ZN(n24946) );
  CKND2D0 U9906 ( .A1(n26976), .A2(n24952), .ZN(n25055) );
  CKND0 U9907 ( .I(n24947), .ZN(n26976) );
  CKND2D0 U9908 ( .A1(n27028), .A2(n27005), .ZN(n24947) );
  OAI222D0 U9909 ( .A1(n25058), .A2(n3947), .B1(n25059), .B2(n3995), .C1(
        n25060), .C2(n3899), .ZN(n27025) );
  CKND2D0 U9910 ( .A1(n26977), .A2(n24952), .ZN(n25058) );
  CKND0 U9911 ( .I(n24944), .ZN(n26977) );
  CKND2D0 U9912 ( .A1(n27006), .A2(n27018), .ZN(n24944) );
  OAI222D0 U9913 ( .A1(n25061), .A2(n4091), .B1(n25062), .B2(n4139), .C1(
        n25063), .C2(n4043), .ZN(n27024) );
  CKND2D0 U9914 ( .A1(n26991), .A2(n24952), .ZN(n25061) );
  NR4D0 U9915 ( .A1(n27029), .A2(n27030), .A3(n27031), .A4(n27032), .ZN(n26962) );
  OAI22D0 U9916 ( .A1(n25068), .A2(n2363), .B1(n25069), .B2(n2891), .ZN(n27032) );
  OAI222D0 U9917 ( .A1(n25070), .A2(n2459), .B1(n25071), .B2(n4283), .C1(
        n25072), .C2(n2603), .ZN(n27031) );
  CKND0 U9918 ( .I(n24937), .ZN(n26981) );
  CKND2D0 U9919 ( .A1(n27004), .A2(n27022), .ZN(n24937) );
  OAI222D0 U9920 ( .A1(n25073), .A2(n4235), .B1(n24930), .B2(n3275), .C1(
        n25074), .C2(n4187), .ZN(n27030) );
  CKND0 U9921 ( .I(n24939), .ZN(n26980) );
  CKND2D0 U9922 ( .A1(n27005), .A2(n27022), .ZN(n24939) );
  NR2D0 U9923 ( .A1(n27019), .A2(n27033), .ZN(n27022) );
  CKND2D0 U9924 ( .A1(n27012), .A2(n27006), .ZN(n24942) );
  NR2D0 U9925 ( .A1(Address[3]), .A2(Address[0]), .ZN(n27006) );
  CKND2D0 U9926 ( .A1(n26982), .A2(n24952), .ZN(n25073) );
  CKND2D0 U9927 ( .A1(n27004), .A2(n27020), .ZN(n24938) );
  OAI222D0 U9928 ( .A1(n24932), .A2(n3371), .B1(n25075), .B2(n4811), .C1(
        n24931), .C2(n3323), .ZN(n27029) );
  CKND2D0 U9929 ( .A1(n27028), .A2(n27012), .ZN(n24941) );
  CKND0 U9930 ( .I(Address[5]), .ZN(n24956) );
  CKND0 U9931 ( .I(Address[6]), .ZN(n24950) );
  NR2D0 U9932 ( .A1(n27023), .A2(Address[5]), .ZN(n26988) );
  CKND0 U9933 ( .I(Address[4]), .ZN(n27023) );
  CKND0 U9934 ( .I(n24943), .ZN(n26998) );
  CKND2D0 U9935 ( .A1(n27028), .A2(n27018), .ZN(n24943) );
  NR2D0 U9936 ( .A1(n27034), .A2(Address[1]), .ZN(n27018) );
  CKND2D0 U9937 ( .A1(n27005), .A2(n27020), .ZN(n24940) );
  NR2D0 U9938 ( .A1(Address[1]), .A2(Address[2]), .ZN(n27005) );
  CKND0 U9939 ( .I(n24936), .ZN(n26983) );
  CKND2D0 U9940 ( .A1(n27012), .A2(n27020), .ZN(n24936) );
  NR2D0 U9941 ( .A1(n27033), .A2(Address[0]), .ZN(n27020) );
  CKND0 U9942 ( .I(Address[3]), .ZN(n27033) );
  NR2D0 U9943 ( .A1(n27035), .A2(n27034), .ZN(n27012) );
  CKND0 U9944 ( .I(Address[2]), .ZN(n27034) );
  CKND0 U9945 ( .I(n24945), .ZN(n26992) );
  CKND2D0 U9946 ( .A1(n27028), .A2(n27004), .ZN(n24945) );
  NR2D0 U9947 ( .A1(n27035), .A2(Address[2]), .ZN(n27004) );
  CKND0 U9948 ( .I(Address[1]), .ZN(n27035) );
  NR2D0 U9949 ( .A1(n27019), .A2(Address[3]), .ZN(n27028) );
  CKND0 U9950 ( .I(Address[0]), .ZN(n27019) );
  CKND0 U9951 ( .I(n24949), .ZN(n24919) );
  NR2D0 U9952 ( .A1(WE), .A2(CS), .ZN(n24949) );
endmodule

