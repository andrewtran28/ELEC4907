
module routing_engine ( port_dest, control, done );
  input [31:0] port_dest;
  output [19:0] control;
  output done;
  wire   \dst[0][1] , \dst[0][0] , \dst[2][2] , \dst[2][1] , \dst[2][0] ,
         \dst[3][2] , \dst[3][0] , \dst[4][2] , \dst[4][1] , \dst[4][0] ,
         \dst[5][2] , \dst[5][1] , \dst[5][0] , \dst[6][2] , \dst[6][1] ,
         \dst[6][0] , \dst[7][1] , \dst[7][0] , N694, N695, N696, N697, N808,
         N810, N811, N922, N923, N924, N925, N1021, N1022, N1023, N1134, N1135,
         N1136, N1137, N1248, N1249, N1250, N1251, N1362, N1363, N1364, N1365,
         N1446, N1447, N1448, \control[13] , n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561;
  assign control[19] = \control[13] ;
  assign control[15] = \control[13] ;
  assign control[13] = \control[13] ;

  LHQD1 \dst_reg[0][1]  ( .E(N694), .D(N696), .Q(\dst[0][1] ) );
  LHQD1 \dst_reg[0][0]  ( .E(N694), .D(N695), .Q(\dst[0][0] ) );
  LHD1 \dst_reg[1][1]  ( .E(N808), .D(N810), .QN(n1561) );
  LHQD1 \dst_reg[2][2]  ( .E(N922), .D(N925), .Q(\dst[2][2] ) );
  LHQD1 \dst_reg[2][1]  ( .E(N922), .D(N924), .Q(\dst[2][1] ) );
  LHQD1 \dst_reg[2][0]  ( .E(N922), .D(N923), .Q(\dst[2][0] ) );
  LHQD1 \dst_reg[3][2]  ( .E(N1021), .D(N1023), .Q(\dst[3][2] ) );
  LHQD1 \dst_reg[3][0]  ( .E(N1021), .D(N1022), .Q(\dst[3][0] ) );
  LHQD1 \dst_reg[4][2]  ( .E(N1134), .D(N1137), .Q(\dst[4][2] ) );
  LHQD1 \dst_reg[4][1]  ( .E(N1134), .D(N1136), .Q(\dst[4][1] ) );
  LHQD1 \dst_reg[4][0]  ( .E(N1134), .D(N1135), .Q(\dst[4][0] ) );
  LHQD1 \dst_reg[5][2]  ( .E(N1248), .D(N1251), .Q(\dst[5][2] ) );
  LHQD1 \dst_reg[5][1]  ( .E(N1248), .D(N1250), .Q(\dst[5][1] ) );
  LHQD1 \dst_reg[5][0]  ( .E(N1248), .D(N1249), .Q(\dst[5][0] ) );
  LHQD1 \dst_reg[6][2]  ( .E(N1362), .D(N1365), .Q(\dst[6][2] ) );
  LHQD1 \dst_reg[6][1]  ( .E(N1362), .D(N1364), .Q(\dst[6][1] ) );
  LHQD1 \dst_reg[6][0]  ( .E(N1362), .D(N1363), .Q(\dst[6][0] ) );
  LHQD1 \dst_reg[7][1]  ( .E(N1446), .D(N1448), .Q(\dst[7][1] ) );
  LHQD1 \dst_reg[7][0]  ( .E(N1446), .D(N1447), .Q(\dst[7][0] ) );
  LHQD2 \dst_reg[1][2]  ( .E(N808), .D(N811), .Q(control[9]) );
  LHQD2 \dst_reg[0][2]  ( .E(N694), .D(N697), .Q(control[11]) );
  MUX2ND2 U868 ( .I0(n1561), .I1(n1191), .S(control[9]), .ZN(control[5]) );
  XOR2D2 U869 ( .A1(n1204), .A2(control[9]), .Z(control[12]) );
  MUX2ND2 U870 ( .I0(n1191), .I1(n1561), .S(control[9]), .ZN(control[4]) );
  MUX3ND0 U871 ( .I0(\dst[6][0] ), .I1(\dst[7][0] ), .I2(n1215), .S0(
        control[16]), .S1(control[14]), .ZN(n1201) );
  XOR2D2 U872 ( .A1(n1216), .A2(control[11]), .Z(control[14]) );
  MUX2ND2 U873 ( .I0(n1195), .I1(n1196), .S(control[7]), .ZN(control[3]) );
  MUX2ND2 U874 ( .I0(n1202), .I1(n1203), .S(control[6]), .ZN(control[1]) );
  CKMUX2D2 U875 ( .I0(n1217), .I1(n1218), .S(\dst[6][2] ), .Z(control[16]) );
  MUX2ND2 U876 ( .I0(n1196), .I1(n1195), .S(control[7]), .ZN(control[2]) );
  IOA21D2 U877 ( .A1(control[11]), .A2(n1197), .B(n1198), .ZN(control[7]) );
  MUX2ND2 U878 ( .I0(n1203), .I1(n1202), .S(control[6]), .ZN(control[0]) );
  CKMUX2D2 U879 ( .I0(\dst[0][1] ), .I1(n1197), .S(n1206), .Z(control[6]) );
  CKMUX2D2 U880 ( .I0(\dst[2][2] ), .I1(\dst[3][2] ), .S(control[18]), .Z(
        control[10]) );
  CKMUX2D2 U881 ( .I0(\dst[3][2] ), .I1(\dst[2][2] ), .S(control[18]), .Z(
        control[8]) );
  AN2D2 U882 ( .A1(n1211), .A2(n1212), .Z(control[18]) );
  MUX4ND2 U883 ( .I0(n1225), .I1(n1226), .I2(n1222), .I3(n1223), .S0(
        \dst[4][1] ), .S1(\dst[4][2] ), .ZN(control[17]) );
  TIEL U884 ( .ZN(\control[13] ) );
  TIEH U885 ( .Z(done) );
  MUX3D0 U886 ( .I0(n1192), .I1(n1193), .I2(n1194), .S0(control[17]), .S1(
        control[12]), .Z(n1191) );
  MUX2ND0 U887 ( .I0(\dst[7][1] ), .I1(\dst[6][1] ), .S(control[16]), .ZN(
        n1194) );
  MUX2ND0 U888 ( .I0(\dst[0][0] ), .I1(n1199), .S(control[11]), .ZN(n1195) );
  MUX2D0 U889 ( .I0(n1200), .I1(n1201), .S(control[10]), .Z(n1196) );
  MUX2ND0 U890 ( .I0(\dst[4][2] ), .I1(\dst[5][2] ), .S(n1205), .ZN(n1204) );
  MUX3ND0 U891 ( .I0(n1192), .I1(n1193), .I2(n1207), .S0(n1205), .S1(
        control[14]), .ZN(n1197) );
  MUX2ND0 U892 ( .I0(\dst[6][1] ), .I1(\dst[7][1] ), .S(control[16]), .ZN(
        n1207) );
  CKND0 U893 ( .I(\dst[4][1] ), .ZN(n1193) );
  CKND0 U894 ( .I(\dst[5][1] ), .ZN(n1192) );
  MUX2ND0 U895 ( .I0(n1199), .I1(\dst[0][0] ), .S(control[11]), .ZN(n1202) );
  MUX3ND0 U896 ( .I0(n1208), .I1(n1209), .I2(n1210), .S0(n1205), .S1(
        control[14]), .ZN(n1199) );
  MUX2ND0 U897 ( .I0(\dst[6][0] ), .I1(\dst[7][0] ), .S(control[16]), .ZN(
        n1210) );
  MUX2D0 U898 ( .I0(n1201), .I1(n1200), .S(control[10]), .Z(n1203) );
  MUX2ND0 U899 ( .I0(\dst[2][0] ), .I1(\dst[3][0] ), .S(control[18]), .ZN(
        n1200) );
  CKXOR2D0 U900 ( .A1(control[11]), .A2(n1213), .Z(n1212) );
  CKXOR2D0 U901 ( .A1(\dst[0][1] ), .A2(n1214), .Z(n1211) );
  MUX2ND0 U902 ( .I0(\dst[5][2] ), .I1(\dst[4][2] ), .S(n1205), .ZN(n1216) );
  OAI21D0 U903 ( .A1(n1219), .A2(n1220), .B(n1221), .ZN(n1218) );
  MUX2D0 U904 ( .I0(n1222), .I1(n1223), .S(\dst[6][1] ), .Z(n1221) );
  CKND0 U905 ( .I(\dst[4][2] ), .ZN(n1219) );
  OAI21D0 U906 ( .A1(\dst[4][2] ), .A2(n1220), .B(n1224), .ZN(n1217) );
  MUX2D0 U907 ( .I0(n1225), .I1(n1226), .S(\dst[6][1] ), .Z(n1224) );
  CKXOR2D0 U908 ( .A1(\dst[6][1] ), .A2(\dst[4][1] ), .Z(n1220) );
  MUX2ND0 U909 ( .I0(n1208), .I1(n1209), .S(n1205), .ZN(n1215) );
  CKND0 U910 ( .I(control[17]), .ZN(n1205) );
  AOI22D0 U911 ( .A1(\dst[2][2] ), .A2(\dst[2][1] ), .B1(control[11]), .B2(
        \dst[0][1] ), .ZN(n1223) );
  AOI22D0 U912 ( .A1(n1214), .A2(\dst[2][2] ), .B1(n1227), .B2(control[11]), 
        .ZN(n1222) );
  OA21D0 U913 ( .A1(\dst[2][2] ), .A2(n1214), .B(n1198), .Z(n1226) );
  CKND2D0 U914 ( .A1(\dst[0][1] ), .A2(n1206), .ZN(n1198) );
  AOI22D0 U915 ( .A1(n1214), .A2(n1213), .B1(n1206), .B2(n1227), .ZN(n1225) );
  CKND0 U916 ( .I(\dst[0][1] ), .ZN(n1227) );
  CKND0 U917 ( .I(control[11]), .ZN(n1206) );
  CKND0 U918 ( .I(\dst[2][2] ), .ZN(n1213) );
  CKND0 U919 ( .I(\dst[2][1] ), .ZN(n1214) );
  CKND0 U920 ( .I(\dst[4][0] ), .ZN(n1209) );
  CKND0 U921 ( .I(\dst[5][0] ), .ZN(n1208) );
  OAI211D0 U922 ( .A1(port_dest[23]), .A2(n1228), .B(n1229), .C(n1230), .ZN(
        N925) );
  AOI21D0 U923 ( .A1(n1231), .A2(port_dest[22]), .B(n1232), .ZN(n1228) );
  OAI221D0 U924 ( .A1(n1233), .A2(n1234), .B1(port_dest[23]), .B2(n1235), .C(
        n1230), .ZN(N924) );
  AOI21D0 U925 ( .A1(n1236), .A2(n1237), .B(n1238), .ZN(n1230) );
  CKND0 U926 ( .I(n1239), .ZN(n1238) );
  NR2D0 U927 ( .A1(n1240), .A2(n1241), .ZN(n1235) );
  AOI21D0 U928 ( .A1(n1242), .A2(n1243), .B(port_dest[23]), .ZN(n1233) );
  CKND2D0 U929 ( .A1(n1244), .A2(n1239), .ZN(N923) );
  ND3D0 U930 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1239) );
  MUX2ND0 U931 ( .I0(n1248), .I1(port_dest[20]), .S(port_dest[23]), .ZN(n1244)
         );
  AOI21D0 U932 ( .A1(n1249), .A2(n1250), .B(n1237), .ZN(n1248) );
  OAI21D0 U933 ( .A1(n1251), .A2(n1240), .B(n1252), .ZN(n1250) );
  INR3D0 U934 ( .A1(n1253), .B1(n1254), .B2(n1255), .ZN(n1240) );
  AOI211D0 U935 ( .A1(n1256), .A2(n1257), .B(n1258), .C(n1241), .ZN(n1251) );
  ND4D0 U936 ( .A1(n1243), .A2(n1255), .A3(n1242), .A4(n1259), .ZN(N922) );
  NR4D0 U937 ( .A1(port_dest[23]), .A2(n1241), .A3(n1237), .A4(n1245), .ZN(
        n1259) );
  CKND0 U938 ( .I(n1260), .ZN(n1245) );
  NR3D0 U939 ( .A1(n1246), .A2(n1261), .A3(n1262), .ZN(n1237) );
  NR2D0 U940 ( .A1(n1253), .A2(n1254), .ZN(n1241) );
  CKND0 U941 ( .I(n1243), .ZN(n1254) );
  CKND0 U942 ( .I(n1232), .ZN(n1242) );
  CKND2D0 U943 ( .A1(n1249), .A2(n1252), .ZN(n1232) );
  CKND2D0 U944 ( .A1(n1263), .A2(n1231), .ZN(n1252) );
  CKND0 U945 ( .I(n1264), .ZN(n1231) );
  CKND2D0 U946 ( .A1(n1261), .A2(n1265), .ZN(n1249) );
  OAI21D0 U947 ( .A1(port_dest[27]), .A2(n1266), .B(n1267), .ZN(N811) );
  AOI221D0 U948 ( .A1(n1268), .A2(n1269), .B1(n1270), .B2(port_dest[26]), .C(
        n1271), .ZN(n1266) );
  OAI222D0 U949 ( .A1(n1272), .A2(n1273), .B1(n1274), .B2(n1275), .C1(n1276), 
        .C2(n1277), .ZN(N810) );
  NR2D0 U950 ( .A1(n1268), .A2(n1278), .ZN(n1274) );
  AOI21D0 U951 ( .A1(n1279), .A2(n1280), .B(port_dest[27]), .ZN(n1272) );
  IND3D0 U952 ( .A1(n1271), .B1(n1281), .B2(n1282), .ZN(N808) );
  CKND0 U953 ( .I(n1268), .ZN(n1282) );
  IOA21D0 U954 ( .A1(n1269), .A2(n1278), .B(n1279), .ZN(n1271) );
  AOI22D0 U955 ( .A1(n1270), .A2(n1283), .B1(n1269), .B2(n1284), .ZN(n1279) );
  CKND0 U956 ( .I(n1285), .ZN(n1270) );
  OAI211D0 U957 ( .A1(port_dest[31]), .A2(n1286), .B(n1287), .C(n1288), .ZN(
        N697) );
  AOI211D0 U958 ( .A1(n1289), .A2(port_dest[30]), .B(n1290), .C(n1291), .ZN(
        n1286) );
  OAI221D0 U959 ( .A1(n1292), .A2(n1293), .B1(port_dest[31]), .B2(n1294), .C(
        n1287), .ZN(N696) );
  OA31D0 U960 ( .A1(n1295), .A2(n1296), .A3(n1290), .B(n1297), .Z(n1292) );
  CKND2D0 U961 ( .A1(n1298), .A2(n1287), .ZN(N695) );
  IND2D0 U962 ( .A1(n1299), .B1(n1300), .ZN(n1287) );
  MUX2ND0 U963 ( .I0(n1301), .I1(port_dest[28]), .S(port_dest[31]), .ZN(n1298)
         );
  NR2D0 U964 ( .A1(n1291), .A2(n1302), .ZN(n1301) );
  MAOI22D0 U965 ( .A1(n1303), .A2(n1304), .B1(n1305), .B2(n1306), .ZN(n1302)
         );
  OAI32D0 U966 ( .A1(n1307), .A2(n1308), .A3(n1295), .B1(n1309), .B2(n1310), 
        .ZN(n1303) );
  NR2D0 U967 ( .A1(n1296), .A2(port_dest[28]), .ZN(n1307) );
  ND4D0 U968 ( .A1(n1299), .A2(n1311), .A3(n1312), .A4(n1313), .ZN(N694) );
  INR2D0 U969 ( .A1(n1294), .B1(n1290), .ZN(n1313) );
  OAI21D0 U970 ( .A1(n1306), .A2(n1305), .B(n1304), .ZN(n1290) );
  IND2D0 U971 ( .A1(n1314), .B1(n1289), .ZN(n1304) );
  AOI211D0 U972 ( .A1(n1315), .A2(n1316), .B(n1308), .C(n1291), .ZN(n1294) );
  INR3D0 U973 ( .A1(n1305), .B1(n1306), .B2(n1317), .ZN(n1291) );
  NR3D0 U974 ( .A1(n1295), .A2(n1296), .A3(n1318), .ZN(n1308) );
  CKND0 U975 ( .I(n1311), .ZN(n1296) );
  CKND2D0 U976 ( .A1(n1319), .A2(n1320), .ZN(N1448) );
  OAI31D0 U977 ( .A1(n1321), .A2(n1322), .A3(n1323), .B(n1324), .ZN(n1320) );
  CKND0 U978 ( .I(n1325), .ZN(n1323) );
  AOI211D0 U979 ( .A1(n1326), .A2(n1327), .B(n1328), .C(n1329), .ZN(n1321) );
  CKND0 U980 ( .I(n1330), .ZN(n1329) );
  CKND2D0 U981 ( .A1(n1331), .A2(port_dest[1]), .ZN(n1327) );
  MUX2ND0 U982 ( .I0(n1332), .I1(n1333), .S(port_dest[3]), .ZN(N1447) );
  AOI21D0 U983 ( .A1(n1334), .A2(n1325), .B(n1322), .ZN(n1332) );
  ND3D0 U984 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1325) );
  OAI21D0 U985 ( .A1(n1328), .A2(n1338), .B(n1330), .ZN(n1334) );
  CKND2D0 U986 ( .A1(n1339), .A2(n1335), .ZN(n1330) );
  AOI32D0 U987 ( .A1(n1340), .A2(n1341), .A3(n1342), .B1(n1343), .B2(n1344), 
        .ZN(n1338) );
  OAI21D0 U988 ( .A1(n1345), .A2(n1346), .B(n1333), .ZN(n1342) );
  ND4D0 U989 ( .A1(n1331), .A2(n1336), .A3(n1326), .A4(n1347), .ZN(N1446) );
  NR4D0 U990 ( .A1(port_dest[3]), .A2(n1328), .A3(n1322), .A4(n1337), .ZN(
        n1347) );
  IINR4D0 U991 ( .A1(n1348), .A2(n1349), .B1(n1337), .B2(n1339), .ZN(n1322) );
  AOI21D0 U992 ( .A1(n1350), .A2(n1351), .B(n1352), .ZN(n1337) );
  INR2D0 U993 ( .A1(n1335), .B1(n1353), .ZN(n1348) );
  AOI211D0 U994 ( .A1(n1354), .A2(n1355), .B(n1343), .C(n1356), .ZN(n1335) );
  CKND0 U995 ( .I(n1357), .ZN(n1343) );
  AN4D0 U996 ( .A1(n1344), .A2(n1355), .A3(n1357), .A4(n1354), .Z(n1328) );
  CKND0 U997 ( .I(n1356), .ZN(n1344) );
  OA21D0 U998 ( .A1(n1356), .A2(n1357), .B(n1340), .Z(n1326) );
  ND3D0 U999 ( .A1(n1358), .A2(n1359), .A3(n1331), .ZN(n1340) );
  OAI21D0 U1000 ( .A1(port_dest[7]), .A2(n1360), .B(n1361), .ZN(n1357) );
  OAI21D0 U1001 ( .A1(n1362), .A2(n1363), .B(n1331), .ZN(n1356) );
  CKND0 U1002 ( .I(n1339), .ZN(n1336) );
  NR2D0 U1003 ( .A1(n1350), .A2(n1351), .ZN(n1339) );
  OA21D0 U1004 ( .A1(n1345), .A2(n1346), .B(n1341), .Z(n1331) );
  CKND2D0 U1005 ( .A1(n1364), .A2(port_dest[7]), .ZN(n1341) );
  OAI221D0 U1006 ( .A1(port_dest[7]), .A2(n1365), .B1(n1366), .B2(n1354), .C(
        n1367), .ZN(N1365) );
  NR2D0 U1007 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
  ND3D0 U1008 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1354) );
  NR2D0 U1009 ( .A1(n1373), .A2(n1374), .ZN(n1365) );
  OAI221D0 U1010 ( .A1(n1375), .A2(n1376), .B1(port_dest[7]), .B2(n1377), .C(
        n1378), .ZN(N1364) );
  AOI21D0 U1011 ( .A1(n1379), .A2(n1380), .B(port_dest[7]), .ZN(n1375) );
  CKND2D0 U1012 ( .A1(n1381), .A2(n1378), .ZN(N1363) );
  CKND0 U1013 ( .I(n1369), .ZN(n1378) );
  NR2D0 U1014 ( .A1(n1349), .A2(n1353), .ZN(n1369) );
  ND3D0 U1015 ( .A1(n1350), .A2(n1352), .A3(n1351), .ZN(n1349) );
  NR2D0 U1016 ( .A1(n1382), .A2(port_dest[7]), .ZN(n1351) );
  MUX2ND0 U1017 ( .I0(n1383), .I1(port_dest[4]), .S(port_dest[7]), .ZN(n1381)
         );
  NR2D0 U1018 ( .A1(n1373), .A2(n1384), .ZN(n1383) );
  AOI22D0 U1019 ( .A1(n1385), .A2(n1386), .B1(n1387), .B2(n1388), .ZN(n1384)
         );
  OAI32D0 U1020 ( .A1(n1389), .A2(n1364), .A3(n1390), .B1(n1360), .B2(n1370), 
        .ZN(n1385) );
  NR2D0 U1021 ( .A1(n1391), .A2(port_dest[4]), .ZN(n1389) );
  ND4D0 U1022 ( .A1(n1362), .A2(n1377), .A3(n1379), .A4(n1353), .ZN(N1362) );
  IND2D0 U1023 ( .A1(n1392), .B1(n1393), .ZN(n1353) );
  CKND0 U1024 ( .I(n1374), .ZN(n1379) );
  OAI21D0 U1025 ( .A1(n1382), .A2(n1350), .B(n1386), .ZN(n1374) );
  ND3D0 U1026 ( .A1(n1372), .A2(n1370), .A3(n1355), .ZN(n1386) );
  CKND0 U1027 ( .I(n1361), .ZN(n1370) );
  CKND0 U1028 ( .I(n1387), .ZN(n1350) );
  AOI211D0 U1029 ( .A1(n1372), .A2(n1361), .B(n1373), .C(n1390), .ZN(n1377) );
  AN2D0 U1030 ( .A1(n1380), .A2(n1358), .Z(n1390) );
  NR3D0 U1031 ( .A1(n1382), .A2(n1387), .A3(n1352), .ZN(n1373) );
  CKND2D0 U1032 ( .A1(n1394), .A2(n1395), .ZN(n1352) );
  AOI21D0 U1033 ( .A1(n1396), .A2(n1397), .B(n1398), .ZN(n1387) );
  CKND0 U1034 ( .I(n1388), .ZN(n1382) );
  NR3D0 U1035 ( .A1(n1361), .A2(n1355), .A3(n1360), .ZN(n1388) );
  NR2D0 U1036 ( .A1(n1396), .A2(n1397), .ZN(n1355) );
  AOI21D0 U1037 ( .A1(n1399), .A2(n1400), .B(n1401), .ZN(n1361) );
  CKND0 U1038 ( .I(n1360), .ZN(n1372) );
  CKND2D0 U1039 ( .A1(n1380), .A2(n1363), .ZN(n1360) );
  CKND0 U1040 ( .I(n1358), .ZN(n1363) );
  NR2D0 U1041 ( .A1(n1402), .A2(n1403), .ZN(n1358) );
  NR2D0 U1042 ( .A1(n1364), .A2(n1391), .ZN(n1380) );
  CKND0 U1043 ( .I(n1359), .ZN(n1362) );
  CKND2D0 U1044 ( .A1(n1345), .A2(n1346), .ZN(n1359) );
  CKND0 U1045 ( .I(n1391), .ZN(n1346) );
  AOI21D0 U1046 ( .A1(n1404), .A2(n1399), .B(n1405), .ZN(n1391) );
  NR2D0 U1047 ( .A1(port_dest[7]), .A2(n1364), .ZN(n1345) );
  NR2D0 U1048 ( .A1(n1404), .A2(n1399), .ZN(n1364) );
  OAI221D0 U1049 ( .A1(n1406), .A2(n1407), .B1(port_dest[11]), .B2(n1408), .C(
        n1409), .ZN(N1251) );
  NR2D0 U1050 ( .A1(n1410), .A2(port_dest[11]), .ZN(n1406) );
  OAI211D0 U1051 ( .A1(port_dest[11]), .A2(n1411), .B(n1412), .C(n1409), .ZN(
        N1250) );
  AOI21D0 U1052 ( .A1(n1413), .A2(n1414), .B(n1415), .ZN(n1411) );
  OAI21D0 U1053 ( .A1(n1416), .A2(n1417), .B(n1418), .ZN(n1414) );
  CKND0 U1054 ( .I(port_dest[9]), .ZN(n1416) );
  CKND2D0 U1055 ( .A1(n1419), .A2(n1409), .ZN(N1249) );
  CKND2D0 U1056 ( .A1(n1392), .A2(n1393), .ZN(n1409) );
  NR2D0 U1057 ( .A1(n1395), .A2(n1394), .ZN(n1392) );
  ND3D0 U1058 ( .A1(n1396), .A2(n1398), .A3(n1397), .ZN(n1395) );
  NR2D0 U1059 ( .A1(n1420), .A2(port_dest[11]), .ZN(n1397) );
  MUX2ND0 U1060 ( .I0(n1421), .I1(port_dest[8]), .S(port_dest[11]), .ZN(n1419)
         );
  AOI21D0 U1061 ( .A1(n1422), .A2(n1423), .B(n1415), .ZN(n1421) );
  OAI22D0 U1062 ( .A1(n1420), .A2(n1396), .B1(n1424), .B2(n1425), .ZN(n1422)
         );
  AOI211D0 U1063 ( .A1(n1405), .A2(n1426), .B(n1427), .C(n1428), .ZN(n1425) );
  CKND0 U1064 ( .I(n1404), .ZN(n1427) );
  IND4D0 U1065 ( .A1(n1393), .B1(n1403), .B2(n1408), .B3(n1418), .ZN(N1248) );
  NR2D0 U1066 ( .A1(n1424), .A2(n1428), .ZN(n1418) );
  NR2D0 U1067 ( .A1(n1402), .A2(n1417), .ZN(n1428) );
  CKND0 U1068 ( .I(n1429), .ZN(n1402) );
  INR2D0 U1069 ( .A1(n1400), .B1(n1401), .ZN(n1424) );
  INR2D0 U1070 ( .A1(n1413), .B1(n1415), .ZN(n1408) );
  AN4D0 U1071 ( .A1(n1394), .A2(n1410), .A3(n1396), .A4(n1398), .Z(n1415) );
  CKND0 U1072 ( .I(n1430), .ZN(n1398) );
  AOI21D0 U1073 ( .A1(n1431), .A2(n1432), .B(n1433), .ZN(n1394) );
  OA21D0 U1074 ( .A1(n1420), .A2(n1396), .B(n1423), .Z(n1413) );
  ND3D0 U1075 ( .A1(n1410), .A2(n1396), .A3(n1430), .ZN(n1423) );
  NR2D0 U1076 ( .A1(n1431), .A2(n1432), .ZN(n1430) );
  CKND0 U1077 ( .I(n1420), .ZN(n1410) );
  OAI21D0 U1078 ( .A1(port_dest[15]), .A2(n1434), .B(n1435), .ZN(n1396) );
  CKND2D0 U1079 ( .A1(n1400), .A2(n1401), .ZN(n1420) );
  AO21D0 U1080 ( .A1(n1436), .A2(n1437), .B(n1438), .Z(n1401) );
  NR2D0 U1081 ( .A1(n1417), .A2(n1429), .ZN(n1400) );
  NR2D0 U1082 ( .A1(n1439), .A2(n1440), .ZN(n1429) );
  NR2D0 U1083 ( .A1(n1417), .A2(port_dest[11]), .ZN(n1403) );
  CKND2D0 U1084 ( .A1(n1404), .A2(n1405), .ZN(n1417) );
  OAI21D0 U1085 ( .A1(port_dest[15]), .A2(n1441), .B(n1442), .ZN(n1405) );
  CKND2D0 U1086 ( .A1(n1441), .A2(port_dest[15]), .ZN(n1404) );
  NR2D0 U1087 ( .A1(n1443), .A2(n1444), .ZN(n1393) );
  OAI211D0 U1088 ( .A1(port_dest[15]), .A2(n1445), .B(n1446), .C(n1447), .ZN(
        N1137) );
  CKND0 U1089 ( .I(n1448), .ZN(n1447) );
  OA21D0 U1090 ( .A1(n1434), .A2(n1449), .B(n1450), .Z(n1445) );
  OAI221D0 U1091 ( .A1(port_dest[15]), .A2(n1451), .B1(n1452), .B2(n1453), .C(
        n1446), .ZN(N1136) );
  MOAI22D0 U1092 ( .A1(port_dest[15]), .A2(n1454), .B1(n1432), .B2(n1455), 
        .ZN(n1453) );
  NR2D0 U1093 ( .A1(n1456), .A2(n1457), .ZN(n1454) );
  INR2D0 U1094 ( .A1(n1458), .B1(n1459), .ZN(n1451) );
  OAI221D0 U1095 ( .A1(n1459), .A2(n1460), .B1(n1436), .B2(n1461), .C(n1446), 
        .ZN(N1135) );
  IND2D0 U1096 ( .A1(n1443), .B1(n1444), .ZN(n1446) );
  AN3D0 U1097 ( .A1(n1433), .A2(n1431), .A3(n1432), .Z(n1444) );
  AOI32D0 U1098 ( .A1(n1462), .A2(n1436), .A3(n1463), .B1(n1455), .B2(n1432), 
        .ZN(n1460) );
  NR2D0 U1099 ( .A1(n1464), .A2(port_dest[15]), .ZN(n1432) );
  OAI32D0 U1100 ( .A1(n1465), .A2(n1441), .A3(n1466), .B1(n1467), .B2(n1438), 
        .ZN(n1463) );
  CKND0 U1101 ( .I(n1468), .ZN(n1441) );
  NR2D0 U1102 ( .A1(n1442), .A2(port_dest[12]), .ZN(n1465) );
  CKND0 U1103 ( .I(n1456), .ZN(n1462) );
  ND4D0 U1104 ( .A1(n1440), .A2(n1458), .A3(n1450), .A4(n1443), .ZN(N1134) );
  OAI31D0 U1105 ( .A1(n1469), .A2(port_dest[19]), .A3(n1470), .B(n1471), .ZN(
        n1443) );
  AOI211D0 U1106 ( .A1(n1472), .A2(n1455), .B(n1456), .C(n1459), .ZN(n1450) );
  NR3D0 U1107 ( .A1(n1464), .A2(n1455), .A3(n1433), .ZN(n1459) );
  OAI21D0 U1108 ( .A1(port_dest[19]), .A2(n1469), .B(n1470), .ZN(n1433) );
  CKND0 U1109 ( .I(n1472), .ZN(n1464) );
  NR2D0 U1110 ( .A1(n1473), .A2(n1434), .ZN(n1456) );
  CKND0 U1111 ( .I(n1431), .ZN(n1455) );
  OAI21D0 U1112 ( .A1(n1474), .A2(n1475), .B(n1476), .ZN(n1431) );
  NR2D0 U1113 ( .A1(n1434), .A2(n1435), .ZN(n1472) );
  CKND0 U1114 ( .I(n1473), .ZN(n1435) );
  CKND2D0 U1115 ( .A1(n1474), .A2(n1475), .ZN(n1473) );
  CKND2D0 U1116 ( .A1(n1437), .A2(n1438), .ZN(n1434) );
  IAO21D0 U1117 ( .A1(n1467), .A2(n1438), .B(n1466), .ZN(n1458) );
  NR2D0 U1118 ( .A1(n1439), .A2(n1457), .ZN(n1466) );
  OAI21D0 U1119 ( .A1(n1477), .A2(n1478), .B(n1479), .ZN(n1438) );
  CKND0 U1120 ( .I(n1437), .ZN(n1467) );
  INR2D0 U1121 ( .A1(n1439), .B1(n1457), .ZN(n1437) );
  CKND2D0 U1122 ( .A1(n1477), .A2(n1478), .ZN(n1439) );
  ND3D0 U1123 ( .A1(n1480), .A2(n1481), .A3(n1482), .ZN(n1478) );
  NR2D0 U1124 ( .A1(n1457), .A2(port_dest[15]), .ZN(n1440) );
  IND2D0 U1125 ( .A1(n1442), .B1(n1468), .ZN(n1457) );
  CKND2D0 U1126 ( .A1(n1483), .A2(port_dest[19]), .ZN(n1468) );
  AOI21D0 U1127 ( .A1(n1480), .A2(n1481), .B(n1482), .ZN(n1442) );
  OAI221D0 U1128 ( .A1(n1484), .A2(n1475), .B1(port_dest[19]), .B2(n1485), .C(
        n1486), .ZN(N1023) );
  CKND0 U1129 ( .I(port_dest[18]), .ZN(n1484) );
  MUX2ND0 U1130 ( .I0(n1487), .I1(n1488), .S(port_dest[19]), .ZN(N1022) );
  INR2D0 U1131 ( .A1(n1489), .B1(n1490), .ZN(n1487) );
  AOI21D0 U1132 ( .A1(n1470), .A2(n1491), .B(n1492), .ZN(n1490) );
  AOI31D0 U1133 ( .A1(n1493), .A2(n1494), .A3(n1476), .B(n1495), .ZN(n1492) );
  AOI221D0 U1134 ( .A1(n1474), .A2(n1493), .B1(n1496), .B2(n1482), .C(n1483), 
        .ZN(n1495) );
  OAI21D0 U1135 ( .A1(port_dest[16]), .A2(n1479), .B(n1497), .ZN(n1496) );
  CKND0 U1136 ( .I(n1477), .ZN(n1497) );
  IND2D0 U1137 ( .A1(n1475), .B1(n1485), .ZN(N1021) );
  AN2D0 U1138 ( .A1(n1489), .A2(n1498), .Z(n1485) );
  OAI31D0 U1139 ( .A1(n1474), .A2(n1470), .A3(n1476), .B(n1493), .ZN(n1498) );
  CKND0 U1140 ( .I(n1499), .ZN(n1476) );
  CKND0 U1141 ( .I(n1494), .ZN(n1474) );
  IND3D0 U1142 ( .A1(n1470), .B1(n1491), .B2(n1471), .ZN(n1489) );
  AOI21D0 U1143 ( .A1(n1246), .A2(n1247), .B(n1260), .ZN(n1471) );
  OAI21D0 U1144 ( .A1(n1278), .A2(n1275), .B(n1268), .ZN(n1260) );
  NR2D0 U1145 ( .A1(n1299), .A2(n1300), .ZN(n1268) );
  INR2D0 U1146 ( .A1(n1317), .B1(n1500), .ZN(n1300) );
  ND4D0 U1147 ( .A1(n1501), .A2(n1502), .A3(n1503), .A4(n1504), .ZN(n1299) );
  AOI33D0 U1148 ( .A1(n1505), .A2(port_dest[10]), .A3(port_dest[8]), .B1(n1506), .B2(port_dest[2]), .B3(port_dest[0]), .ZN(n1504) );
  AOI33D0 U1149 ( .A1(port_dest[12]), .A2(n1448), .A3(port_dest[13]), .B1(
        port_dest[16]), .B2(n1507), .B3(port_dest[17]), .ZN(n1503) );
  AOI33D0 U1150 ( .A1(port_dest[4]), .A2(n1368), .A3(port_dest[5]), .B1(
        port_dest[28]), .B2(n1508), .B3(port_dest[29]), .ZN(n1502) );
  AOI33D0 U1151 ( .A1(port_dest[20]), .A2(n1509), .A3(port_dest[21]), .B1(
        port_dest[24]), .B2(n1510), .B3(port_dest[25]), .ZN(n1501) );
  CKND0 U1152 ( .I(n1469), .ZN(n1491) );
  ND3D0 U1153 ( .A1(n1494), .A2(n1499), .A3(n1493), .ZN(n1469) );
  OAI21D0 U1154 ( .A1(port_dest[23]), .A2(n1262), .B(n1261), .ZN(n1499) );
  OAI21D0 U1155 ( .A1(port_dest[23]), .A2(n1264), .B(n1263), .ZN(n1494) );
  NR2D0 U1156 ( .A1(n1246), .A2(n1247), .ZN(n1470) );
  NR3D0 U1157 ( .A1(n1261), .A2(port_dest[23]), .A3(n1262), .ZN(n1247) );
  CKND0 U1158 ( .I(n1265), .ZN(n1262) );
  NR2D0 U1159 ( .A1(n1264), .A2(n1263), .ZN(n1265) );
  INR2D0 U1160 ( .A1(n1283), .B1(n1281), .ZN(n1263) );
  NR2D0 U1161 ( .A1(n1285), .A2(port_dest[27]), .ZN(n1281) );
  ND3D0 U1162 ( .A1(n1255), .A2(n1253), .A3(n1243), .ZN(n1264) );
  AOI21D0 U1163 ( .A1(n1511), .A2(n1269), .B(n1512), .ZN(n1261) );
  CKND2D0 U1164 ( .A1(n1278), .A2(n1275), .ZN(n1246) );
  ND3D0 U1165 ( .A1(n1512), .A2(n1511), .A3(n1269), .ZN(n1275) );
  NR2D0 U1166 ( .A1(n1285), .A2(n1283), .ZN(n1269) );
  AOI21D0 U1167 ( .A1(n1297), .A2(n1289), .B(n1314), .ZN(n1283) );
  CKND2D0 U1168 ( .A1(n1280), .A2(n1276), .ZN(n1285) );
  NR2D0 U1169 ( .A1(n1513), .A2(n1514), .ZN(n1276) );
  CKND0 U1170 ( .I(n1284), .ZN(n1512) );
  NR2D0 U1171 ( .A1(n1305), .A2(n1515), .ZN(n1284) );
  INR2D0 U1172 ( .A1(n1500), .B1(n1317), .ZN(n1278) );
  ND4D0 U1173 ( .A1(n1516), .A2(n1517), .A3(n1518), .A4(n1519), .ZN(n1317) );
  AOI33D0 U1174 ( .A1(port_dest[10]), .A2(n1426), .A3(n1505), .B1(port_dest[2]), .B2(n1333), .B3(n1506), .ZN(n1519) );
  AOI33D0 U1175 ( .A1(n1448), .A2(n1461), .A3(port_dest[13]), .B1(n1507), .B2(
        n1488), .B3(port_dest[17]), .ZN(n1518) );
  AOI33D0 U1176 ( .A1(n1368), .A2(n1520), .A3(port_dest[5]), .B1(n1508), .B2(
        n1521), .B3(port_dest[29]), .ZN(n1517) );
  AOI33D0 U1177 ( .A1(n1509), .A2(n1256), .A3(port_dest[21]), .B1(n1510), .B2(
        n1522), .B3(port_dest[25]), .ZN(n1516) );
  CKND2D0 U1178 ( .A1(n1515), .A2(n1305), .ZN(n1500) );
  ND4D0 U1179 ( .A1(n1523), .A2(n1524), .A3(n1525), .A4(n1526), .ZN(n1305) );
  AOI33D0 U1180 ( .A1(port_dest[10]), .A2(n1527), .A3(port_dest[8]), .B1(
        port_dest[2]), .B2(n1528), .B3(port_dest[0]), .ZN(n1526) );
  AOI33D0 U1181 ( .A1(n1448), .A2(n1452), .A3(port_dest[12]), .B1(n1507), .B2(
        n1529), .B3(port_dest[16]), .ZN(n1525) );
  AOI33D0 U1182 ( .A1(n1368), .A2(n1376), .A3(port_dest[4]), .B1(n1508), .B2(
        n1293), .B3(port_dest[28]), .ZN(n1524) );
  AOI33D0 U1183 ( .A1(n1509), .A2(n1234), .A3(port_dest[20]), .B1(n1510), .B2(
        n1273), .B3(port_dest[24]), .ZN(n1523) );
  NR2D0 U1184 ( .A1(n1306), .A2(port_dest[31]), .ZN(n1515) );
  CKND2D0 U1185 ( .A1(n1289), .A2(n1314), .ZN(n1306) );
  ND4D0 U1186 ( .A1(n1530), .A2(n1531), .A3(n1532), .A4(n1533), .ZN(n1314) );
  AOI33D0 U1187 ( .A1(n1527), .A2(n1426), .A3(port_dest[10]), .B1(n1528), .B2(
        n1333), .B3(port_dest[2]), .ZN(n1533) );
  AOI33D0 U1188 ( .A1(n1461), .A2(n1452), .A3(n1448), .B1(n1488), .B2(n1529), 
        .B3(n1507), .ZN(n1532) );
  CKND0 U1189 ( .I(n1486), .ZN(n1507) );
  CKND2D0 U1190 ( .A1(port_dest[19]), .A2(port_dest[18]), .ZN(n1486) );
  NR2D0 U1191 ( .A1(n1436), .A2(n1449), .ZN(n1448) );
  CKND0 U1192 ( .I(port_dest[14]), .ZN(n1449) );
  AOI33D0 U1193 ( .A1(n1520), .A2(n1376), .A3(n1368), .B1(n1521), .B2(n1293), 
        .B3(n1508), .ZN(n1531) );
  CKND0 U1194 ( .I(n1288), .ZN(n1508) );
  CKND2D0 U1195 ( .A1(port_dest[31]), .A2(port_dest[30]), .ZN(n1288) );
  NR2D0 U1196 ( .A1(n1371), .A2(n1366), .ZN(n1368) );
  CKND0 U1197 ( .I(port_dest[6]), .ZN(n1366) );
  AOI33D0 U1198 ( .A1(n1256), .A2(n1234), .A3(n1509), .B1(n1522), .B2(n1273), 
        .B3(n1510), .ZN(n1530) );
  CKND0 U1199 ( .I(n1267), .ZN(n1510) );
  CKND2D0 U1200 ( .A1(port_dest[27]), .A2(port_dest[26]), .ZN(n1267) );
  CKND0 U1201 ( .I(n1229), .ZN(n1509) );
  CKND2D0 U1202 ( .A1(port_dest[23]), .A2(port_dest[22]), .ZN(n1229) );
  NR2D0 U1203 ( .A1(n1309), .A2(n1316), .ZN(n1289) );
  CKND0 U1204 ( .I(n1310), .ZN(n1316) );
  CKND2D0 U1205 ( .A1(n1493), .A2(n1481), .ZN(n1475) );
  INR4D0 U1206 ( .A1(n1482), .B1(n1479), .B2(n1483), .B3(n1477), .ZN(n1493) );
  AOI21D0 U1207 ( .A1(n1236), .A2(n1243), .B(n1253), .ZN(n1477) );
  CKND0 U1208 ( .I(n1480), .ZN(n1483) );
  CKND2D0 U1209 ( .A1(n1258), .A2(port_dest[23]), .ZN(n1480) );
  AOI31D0 U1210 ( .A1(n1243), .A2(n1236), .A3(n1253), .B(n1255), .ZN(n1479) );
  OAI21D0 U1211 ( .A1(n1514), .A2(n1277), .B(n1513), .ZN(n1255) );
  AOI21D0 U1212 ( .A1(n1297), .A2(n1315), .B(n1310), .ZN(n1513) );
  ND4D0 U1213 ( .A1(n1534), .A2(n1535), .A3(n1536), .A4(n1537), .ZN(n1310) );
  AOI33D0 U1214 ( .A1(port_dest[16]), .A2(n1538), .A3(port_dest[17]), .B1(
        port_dest[12]), .B2(n1539), .B3(port_dest[13]), .ZN(n1537) );
  AOI33D0 U1215 ( .A1(port_dest[4]), .A2(n1540), .A3(port_dest[5]), .B1(
        port_dest[24]), .B2(n1541), .B3(port_dest[25]), .ZN(n1536) );
  AOI33D0 U1216 ( .A1(port_dest[28]), .A2(n1542), .A3(port_dest[29]), .B1(
        port_dest[20]), .B2(n1543), .B3(port_dest[21]), .ZN(n1535) );
  AOI33D0 U1217 ( .A1(n1505), .A2(n1407), .A3(port_dest[8]), .B1(n1506), .B2(
        n1544), .B3(port_dest[0]), .ZN(n1534) );
  CKND0 U1218 ( .I(n1309), .ZN(n1315) );
  ND3D0 U1219 ( .A1(n1545), .A2(n1311), .A3(n1318), .ZN(n1309) );
  CKND2D0 U1220 ( .A1(n1514), .A2(n1277), .ZN(n1253) );
  CKND2D0 U1221 ( .A1(n1280), .A2(n1511), .ZN(n1277) );
  AOI21D0 U1222 ( .A1(port_dest[31]), .A2(n1295), .B(n1546), .ZN(n1280) );
  AOI21D0 U1223 ( .A1(n1311), .A2(n1312), .B(n1318), .ZN(n1514) );
  ND4D0 U1224 ( .A1(n1547), .A2(n1548), .A3(n1549), .A4(n1550), .ZN(n1318) );
  AOI33D0 U1225 ( .A1(n1538), .A2(n1488), .A3(port_dest[17]), .B1(n1539), .B2(
        n1461), .B3(port_dest[13]), .ZN(n1550) );
  AOI33D0 U1226 ( .A1(n1540), .A2(n1520), .A3(port_dest[5]), .B1(n1541), .B2(
        n1522), .B3(port_dest[25]), .ZN(n1549) );
  AOI33D0 U1227 ( .A1(n1542), .A2(n1521), .A3(port_dest[29]), .B1(n1543), .B2(
        n1256), .B3(port_dest[21]), .ZN(n1548) );
  AOI33D0 U1228 ( .A1(n1407), .A2(n1426), .A3(n1505), .B1(n1333), .B2(n1544), 
        .B3(n1506), .ZN(n1547) );
  CKND0 U1229 ( .I(n1319), .ZN(n1506) );
  CKND2D0 U1230 ( .A1(port_dest[1]), .A2(port_dest[3]), .ZN(n1319) );
  CKND0 U1231 ( .I(n1412), .ZN(n1505) );
  CKND2D0 U1232 ( .A1(port_dest[9]), .A2(port_dest[11]), .ZN(n1412) );
  NR2D0 U1233 ( .A1(n1258), .A2(n1551), .ZN(n1243) );
  OAI21D0 U1234 ( .A1(port_dest[23]), .A2(n1258), .B(n1551), .ZN(n1482) );
  CKND0 U1235 ( .I(n1257), .ZN(n1551) );
  OAI21D0 U1236 ( .A1(n1552), .A2(port_dest[27]), .B(n1546), .ZN(n1257) );
  NR2D0 U1237 ( .A1(n1311), .A2(n1312), .ZN(n1546) );
  NR2D0 U1238 ( .A1(port_dest[31]), .A2(n1295), .ZN(n1312) );
  CKND0 U1239 ( .I(n1545), .ZN(n1295) );
  ND4D0 U1240 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .ZN(n1311) );
  AOI33D0 U1241 ( .A1(n1538), .A2(n1529), .A3(port_dest[16]), .B1(n1539), .B2(
        n1452), .B3(port_dest[12]), .ZN(n1556) );
  AOI33D0 U1242 ( .A1(n1527), .A2(n1407), .A3(port_dest[8]), .B1(n1540), .B2(
        n1376), .B3(port_dest[4]), .ZN(n1555) );
  AOI33D0 U1243 ( .A1(n1528), .A2(n1544), .A3(port_dest[0]), .B1(n1541), .B2(
        n1273), .B3(port_dest[24]), .ZN(n1554) );
  AOI33D0 U1244 ( .A1(n1542), .A2(n1293), .A3(port_dest[28]), .B1(n1543), .B2(
        n1234), .B3(port_dest[20]), .ZN(n1553) );
  NR2D0 U1245 ( .A1(n1297), .A2(n1545), .ZN(n1552) );
  NR3D0 U1246 ( .A1(n1511), .A2(n1297), .A3(n1545), .ZN(n1258) );
  ND4D0 U1247 ( .A1(n1557), .A2(n1558), .A3(n1559), .A4(n1560), .ZN(n1545) );
  AOI33D0 U1248 ( .A1(n1488), .A2(n1529), .A3(n1538), .B1(n1461), .B2(n1452), 
        .B3(n1539), .ZN(n1560) );
  NR2D0 U1249 ( .A1(n1436), .A2(port_dest[14]), .ZN(n1539) );
  CKND0 U1250 ( .I(port_dest[15]), .ZN(n1436) );
  CKND0 U1251 ( .I(port_dest[13]), .ZN(n1452) );
  CKND0 U1252 ( .I(port_dest[12]), .ZN(n1461) );
  NR2D0 U1253 ( .A1(n1481), .A2(port_dest[18]), .ZN(n1538) );
  CKND0 U1254 ( .I(port_dest[19]), .ZN(n1481) );
  CKND0 U1255 ( .I(port_dest[17]), .ZN(n1529) );
  CKND0 U1256 ( .I(port_dest[16]), .ZN(n1488) );
  AOI33D0 U1257 ( .A1(n1407), .A2(n1426), .A3(n1527), .B1(n1520), .B2(n1376), 
        .B3(n1540), .ZN(n1559) );
  NR2D0 U1258 ( .A1(n1371), .A2(port_dest[6]), .ZN(n1540) );
  CKND0 U1259 ( .I(port_dest[7]), .ZN(n1371) );
  CKND0 U1260 ( .I(port_dest[5]), .ZN(n1376) );
  CKND0 U1261 ( .I(port_dest[4]), .ZN(n1520) );
  NR2D0 U1262 ( .A1(n1399), .A2(port_dest[9]), .ZN(n1527) );
  CKND0 U1263 ( .I(port_dest[11]), .ZN(n1399) );
  CKND0 U1264 ( .I(port_dest[8]), .ZN(n1426) );
  CKND0 U1265 ( .I(port_dest[10]), .ZN(n1407) );
  AOI33D0 U1266 ( .A1(n1333), .A2(n1544), .A3(n1528), .B1(n1522), .B2(n1273), 
        .B3(n1541), .ZN(n1558) );
  NR2D0 U1267 ( .A1(n1511), .A2(port_dest[26]), .ZN(n1541) );
  CKND0 U1268 ( .I(port_dest[25]), .ZN(n1273) );
  CKND0 U1269 ( .I(port_dest[24]), .ZN(n1522) );
  NR2D0 U1270 ( .A1(n1324), .A2(port_dest[1]), .ZN(n1528) );
  CKND0 U1271 ( .I(port_dest[3]), .ZN(n1324) );
  CKND0 U1272 ( .I(port_dest[2]), .ZN(n1544) );
  CKND0 U1273 ( .I(port_dest[0]), .ZN(n1333) );
  AOI33D0 U1274 ( .A1(n1521), .A2(n1293), .A3(n1542), .B1(n1256), .B2(n1234), 
        .B3(n1543), .ZN(n1557) );
  NR2D0 U1275 ( .A1(n1236), .A2(port_dest[22]), .ZN(n1543) );
  CKND0 U1276 ( .I(port_dest[23]), .ZN(n1236) );
  CKND0 U1277 ( .I(port_dest[21]), .ZN(n1234) );
  CKND0 U1278 ( .I(port_dest[20]), .ZN(n1256) );
  NR2D0 U1279 ( .A1(n1297), .A2(port_dest[30]), .ZN(n1542) );
  CKND0 U1280 ( .I(port_dest[29]), .ZN(n1293) );
  CKND0 U1281 ( .I(port_dest[28]), .ZN(n1521) );
  CKND0 U1282 ( .I(port_dest[31]), .ZN(n1297) );
  CKND0 U1283 ( .I(port_dest[27]), .ZN(n1511) );
endmodule

