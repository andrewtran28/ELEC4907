
module routingCache ( clk, rst, wr, val, tag, vld, cfg );
  input [19:0] val;
  input [23:0] tag;
  output [19:0] cfg;
  input clk, rst, wr;
  output vld;
  wire   \entry[7][43] , \entry[7][42] , \entry[7][41] , \entry[7][40] ,
         \entry[7][39] , \entry[7][38] , \entry[7][37] , \entry[7][36] ,
         \entry[7][35] , \entry[7][34] , \entry[7][33] , \entry[7][32] ,
         \entry[7][31] , \entry[7][30] , \entry[7][29] , \entry[7][28] ,
         \entry[7][27] , \entry[7][26] , \entry[7][25] , \entry[7][24] ,
         \entry[7][23] , \entry[7][22] , \entry[7][21] , \entry[7][20] ,
         \entry[7][19] , \entry[7][18] , \entry[7][17] , \entry[7][16] ,
         \entry[7][15] , \entry[7][14] , \entry[7][13] , \entry[7][12] ,
         \entry[7][11] , \entry[7][10] , \entry[7][9] , \entry[7][8] ,
         \entry[7][7] , \entry[7][6] , \entry[7][5] , \entry[7][4] ,
         \entry[7][3] , \entry[7][2] , \entry[7][1] , \entry[7][0] ,
         \entry[6][43] , \entry[6][42] , \entry[6][41] , \entry[6][40] ,
         \entry[6][39] , \entry[6][38] , \entry[6][37] , \entry[6][36] ,
         \entry[6][35] , \entry[6][34] , \entry[6][33] , \entry[6][32] ,
         \entry[6][31] , \entry[6][30] , \entry[6][29] , \entry[6][28] ,
         \entry[6][27] , \entry[6][26] , \entry[6][25] , \entry[6][24] ,
         \entry[6][23] , \entry[6][22] , \entry[6][21] , \entry[6][20] ,
         \entry[6][19] , \entry[6][18] , \entry[6][17] , \entry[6][16] ,
         \entry[6][15] , \entry[6][14] , \entry[6][13] , \entry[6][12] ,
         \entry[6][11] , \entry[6][10] , \entry[6][9] , \entry[6][8] ,
         \entry[6][7] , \entry[6][6] , \entry[6][5] , \entry[6][4] ,
         \entry[6][3] , \entry[6][2] , \entry[6][1] , \entry[6][0] ,
         \entry[5][43] , \entry[5][42] , \entry[5][41] , \entry[5][40] ,
         \entry[5][39] , \entry[5][38] , \entry[5][37] , \entry[5][36] ,
         \entry[5][35] , \entry[5][34] , \entry[5][33] , \entry[5][32] ,
         \entry[5][31] , \entry[5][30] , \entry[5][29] , \entry[5][28] ,
         \entry[5][27] , \entry[5][26] , \entry[5][25] , \entry[5][24] ,
         \entry[5][23] , \entry[5][22] , \entry[5][21] , \entry[5][20] ,
         \entry[5][19] , \entry[5][18] , \entry[5][17] , \entry[5][16] ,
         \entry[5][15] , \entry[5][14] , \entry[5][13] , \entry[5][12] ,
         \entry[5][11] , \entry[5][10] , \entry[5][9] , \entry[5][8] ,
         \entry[5][7] , \entry[5][6] , \entry[5][5] , \entry[5][4] ,
         \entry[5][3] , \entry[5][2] , \entry[5][1] , \entry[5][0] ,
         \entry[4][43] , \entry[4][42] , \entry[4][41] , \entry[4][40] ,
         \entry[4][39] , \entry[4][38] , \entry[4][37] , \entry[4][36] ,
         \entry[4][35] , \entry[4][34] , \entry[4][33] , \entry[4][32] ,
         \entry[4][31] , \entry[4][30] , \entry[4][29] , \entry[4][28] ,
         \entry[4][27] , \entry[4][26] , \entry[4][25] , \entry[4][24] ,
         \entry[4][23] , \entry[4][22] , \entry[4][21] , \entry[4][20] ,
         \entry[4][19] , \entry[4][18] , \entry[4][17] , \entry[4][16] ,
         \entry[4][15] , \entry[4][14] , \entry[4][13] , \entry[4][12] ,
         \entry[4][11] , \entry[4][10] , \entry[4][9] , \entry[4][8] ,
         \entry[4][7] , \entry[4][6] , \entry[4][5] , \entry[4][4] ,
         \entry[4][3] , \entry[4][2] , \entry[4][1] , \entry[4][0] ,
         \entry[3][43] , \entry[3][42] , \entry[3][41] , \entry[3][40] ,
         \entry[3][39] , \entry[3][38] , \entry[3][37] , \entry[3][36] ,
         \entry[3][35] , \entry[3][34] , \entry[3][33] , \entry[3][32] ,
         \entry[3][31] , \entry[3][30] , \entry[3][29] , \entry[3][28] ,
         \entry[3][27] , \entry[3][26] , \entry[3][25] , \entry[3][24] ,
         \entry[3][23] , \entry[3][22] , \entry[3][21] , \entry[3][20] ,
         \entry[3][19] , \entry[3][18] , \entry[3][17] , \entry[3][16] ,
         \entry[3][15] , \entry[3][14] , \entry[3][13] , \entry[3][12] ,
         \entry[3][11] , \entry[3][10] , \entry[3][9] , \entry[3][8] ,
         \entry[3][7] , \entry[3][6] , \entry[3][5] , \entry[3][4] ,
         \entry[3][3] , \entry[3][2] , \entry[3][1] , \entry[3][0] ,
         \entry[2][43] , \entry[2][42] , \entry[2][41] , \entry[2][40] ,
         \entry[2][39] , \entry[2][38] , \entry[2][37] , \entry[2][36] ,
         \entry[2][35] , \entry[2][34] , \entry[2][33] , \entry[2][32] ,
         \entry[2][31] , \entry[2][30] , \entry[2][29] , \entry[2][28] ,
         \entry[2][27] , \entry[2][26] , \entry[2][25] , \entry[2][24] ,
         \entry[2][23] , \entry[2][22] , \entry[2][21] , \entry[2][20] ,
         \entry[2][19] , \entry[2][18] , \entry[2][17] , \entry[2][16] ,
         \entry[2][15] , \entry[2][14] , \entry[2][13] , \entry[2][12] ,
         \entry[2][11] , \entry[2][10] , \entry[2][9] , \entry[2][8] ,
         \entry[2][7] , \entry[2][6] , \entry[2][5] , \entry[2][4] ,
         \entry[2][3] , \entry[2][2] , \entry[2][1] , \entry[2][0] ,
         \entry[1][43] , \entry[1][42] , \entry[1][41] , \entry[1][40] ,
         \entry[1][39] , \entry[1][38] , \entry[1][37] , \entry[1][36] ,
         \entry[1][35] , \entry[1][34] , \entry[1][33] , \entry[1][32] ,
         \entry[1][31] , \entry[1][30] , \entry[1][29] , \entry[1][28] ,
         \entry[1][27] , \entry[1][26] , \entry[1][25] , \entry[1][24] ,
         \entry[1][23] , \entry[1][22] , \entry[1][21] , \entry[1][20] ,
         \entry[1][19] , \entry[1][18] , \entry[1][17] , \entry[1][16] ,
         \entry[1][15] , \entry[1][14] , \entry[1][13] , \entry[1][12] ,
         \entry[1][11] , \entry[1][10] , \entry[1][9] , \entry[1][8] ,
         \entry[1][7] , \entry[1][6] , \entry[1][5] , \entry[1][4] ,
         \entry[1][3] , \entry[1][2] , \entry[1][1] , \entry[1][0] ,
         \entry[0][43] , \entry[0][42] , \entry[0][41] , \entry[0][40] ,
         \entry[0][39] , \entry[0][38] , \entry[0][37] , \entry[0][36] ,
         \entry[0][35] , \entry[0][34] , \entry[0][33] , \entry[0][32] ,
         \entry[0][31] , \entry[0][30] , \entry[0][29] , \entry[0][28] ,
         \entry[0][27] , \entry[0][26] , \entry[0][25] , \entry[0][24] ,
         \entry[0][23] , \entry[0][22] , \entry[0][21] , \entry[0][20] ,
         \entry[0][19] , \entry[0][18] , \entry[0][17] , \entry[0][16] ,
         \entry[0][15] , \entry[0][14] , \entry[0][13] , \entry[0][12] ,
         \entry[0][11] , \entry[0][10] , \entry[0][9] , \entry[0][8] ,
         \entry[0][7] , \entry[0][6] , \entry[0][5] , \entry[0][4] ,
         \entry[0][3] , \entry[0][2] , \entry[0][1] , \entry[0][0] , N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780;
  wire   [2:0] count;

  EDFQD2 \cfg_reg[19]  ( .D(N125), .E(N105), .CP(clk), .Q(cfg[19]) );
  EDFQD2 \cfg_reg[18]  ( .D(N124), .E(N105), .CP(clk), .Q(cfg[18]) );
  EDFQD2 \cfg_reg[17]  ( .D(N123), .E(N105), .CP(clk), .Q(cfg[17]) );
  EDFQD2 \cfg_reg[16]  ( .D(N122), .E(N105), .CP(clk), .Q(cfg[16]) );
  EDFQD2 \cfg_reg[15]  ( .D(N121), .E(N105), .CP(clk), .Q(cfg[15]) );
  EDFQD2 \cfg_reg[14]  ( .D(N120), .E(N105), .CP(clk), .Q(cfg[14]) );
  EDFQD2 \cfg_reg[13]  ( .D(N119), .E(N105), .CP(clk), .Q(cfg[13]) );
  EDFQD2 \cfg_reg[12]  ( .D(N118), .E(N105), .CP(clk), .Q(cfg[12]) );
  EDFQD2 \cfg_reg[11]  ( .D(N117), .E(N105), .CP(clk), .Q(cfg[11]) );
  EDFQD2 \cfg_reg[10]  ( .D(N116), .E(N105), .CP(clk), .Q(cfg[10]) );
  EDFQD2 \cfg_reg[9]  ( .D(N115), .E(N105), .CP(clk), .Q(cfg[9]) );
  EDFQD2 \cfg_reg[8]  ( .D(N114), .E(N105), .CP(clk), .Q(cfg[8]) );
  EDFQD2 \cfg_reg[7]  ( .D(N113), .E(N105), .CP(clk), .Q(cfg[7]) );
  EDFQD2 \cfg_reg[6]  ( .D(N112), .E(N105), .CP(clk), .Q(cfg[6]) );
  EDFQD2 \cfg_reg[5]  ( .D(N111), .E(N105), .CP(clk), .Q(cfg[5]) );
  EDFQD2 \cfg_reg[4]  ( .D(N110), .E(N105), .CP(clk), .Q(cfg[4]) );
  EDFQD2 \cfg_reg[3]  ( .D(N109), .E(N105), .CP(clk), .Q(cfg[3]) );
  EDFQD2 \cfg_reg[2]  ( .D(N108), .E(N105), .CP(clk), .Q(cfg[2]) );
  EDFQD2 \cfg_reg[1]  ( .D(N107), .E(N105), .CP(clk), .Q(cfg[1]) );
  EDFQD2 \cfg_reg[0]  ( .D(N106), .E(N105), .CP(clk), .Q(cfg[0]) );
  EDFQD1 \count_reg[0]  ( .D(N102), .E(N101), .CP(clk), .Q(count[0]) );
  EDFQD1 \count_reg[1]  ( .D(N103), .E(N101), .CP(clk), .Q(count[1]) );
  EDFQD1 \count_reg[2]  ( .D(N104), .E(N101), .CP(clk), .Q(count[2]) );
  EDFQD1 \entry_reg[7][43]  ( .D(N93), .E(N100), .CP(clk), .Q(\entry[7][43] )
         );
  EDFQD1 \entry_reg[7][42]  ( .D(N92), .E(N100), .CP(clk), .Q(\entry[7][42] )
         );
  EDFQD1 \entry_reg[7][41]  ( .D(N91), .E(N100), .CP(clk), .Q(\entry[7][41] )
         );
  EDFQD1 \entry_reg[7][40]  ( .D(N90), .E(N100), .CP(clk), .Q(\entry[7][40] )
         );
  EDFQD1 \entry_reg[7][39]  ( .D(N89), .E(N100), .CP(clk), .Q(\entry[7][39] )
         );
  EDFQD1 \entry_reg[7][38]  ( .D(N88), .E(N100), .CP(clk), .Q(\entry[7][38] )
         );
  EDFQD1 \entry_reg[7][37]  ( .D(N87), .E(N100), .CP(clk), .Q(\entry[7][37] )
         );
  EDFQD1 \entry_reg[7][36]  ( .D(N86), .E(N100), .CP(clk), .Q(\entry[7][36] )
         );
  EDFQD1 \entry_reg[7][35]  ( .D(N85), .E(N100), .CP(clk), .Q(\entry[7][35] )
         );
  EDFQD1 \entry_reg[7][34]  ( .D(N84), .E(N100), .CP(clk), .Q(\entry[7][34] )
         );
  EDFQD1 \entry_reg[7][33]  ( .D(N83), .E(N100), .CP(clk), .Q(\entry[7][33] )
         );
  EDFQD1 \entry_reg[7][32]  ( .D(N82), .E(N100), .CP(clk), .Q(\entry[7][32] )
         );
  EDFQD1 \entry_reg[7][31]  ( .D(N81), .E(N100), .CP(clk), .Q(\entry[7][31] )
         );
  EDFQD1 \entry_reg[7][30]  ( .D(N80), .E(N100), .CP(clk), .Q(\entry[7][30] )
         );
  EDFQD1 \entry_reg[7][29]  ( .D(N79), .E(N100), .CP(clk), .Q(\entry[7][29] )
         );
  EDFQD1 \entry_reg[7][28]  ( .D(N78), .E(N100), .CP(clk), .Q(\entry[7][28] )
         );
  EDFQD1 \entry_reg[7][27]  ( .D(N77), .E(N100), .CP(clk), .Q(\entry[7][27] )
         );
  EDFQD1 \entry_reg[7][26]  ( .D(N76), .E(N100), .CP(clk), .Q(\entry[7][26] )
         );
  EDFQD1 \entry_reg[7][25]  ( .D(N75), .E(N100), .CP(clk), .Q(\entry[7][25] )
         );
  EDFQD1 \entry_reg[7][24]  ( .D(N74), .E(N100), .CP(clk), .Q(\entry[7][24] )
         );
  EDFQD1 \entry_reg[7][23]  ( .D(N73), .E(N100), .CP(clk), .Q(\entry[7][23] )
         );
  EDFQD1 \entry_reg[7][22]  ( .D(N72), .E(N100), .CP(clk), .Q(\entry[7][22] )
         );
  EDFQD1 \entry_reg[7][21]  ( .D(N71), .E(N100), .CP(clk), .Q(\entry[7][21] )
         );
  EDFQD1 \entry_reg[7][20]  ( .D(N70), .E(N100), .CP(clk), .Q(\entry[7][20] )
         );
  EDFQD1 \entry_reg[7][19]  ( .D(N69), .E(N100), .CP(clk), .Q(\entry[7][19] )
         );
  EDFQD1 \entry_reg[7][18]  ( .D(N68), .E(N100), .CP(clk), .Q(\entry[7][18] )
         );
  EDFQD1 \entry_reg[7][17]  ( .D(N67), .E(N100), .CP(clk), .Q(\entry[7][17] )
         );
  EDFQD1 \entry_reg[7][16]  ( .D(N66), .E(N100), .CP(clk), .Q(\entry[7][16] )
         );
  EDFQD1 \entry_reg[7][15]  ( .D(N65), .E(N100), .CP(clk), .Q(\entry[7][15] )
         );
  EDFQD1 \entry_reg[7][14]  ( .D(N64), .E(N100), .CP(clk), .Q(\entry[7][14] )
         );
  EDFQD1 \entry_reg[7][13]  ( .D(N63), .E(N100), .CP(clk), .Q(\entry[7][13] )
         );
  EDFQD1 \entry_reg[7][12]  ( .D(N62), .E(N100), .CP(clk), .Q(\entry[7][12] )
         );
  EDFQD1 \entry_reg[7][11]  ( .D(N61), .E(N100), .CP(clk), .Q(\entry[7][11] )
         );
  EDFQD1 \entry_reg[7][10]  ( .D(N60), .E(N100), .CP(clk), .Q(\entry[7][10] )
         );
  EDFQD1 \entry_reg[7][9]  ( .D(N59), .E(N100), .CP(clk), .Q(\entry[7][9] ) );
  EDFQD1 \entry_reg[7][8]  ( .D(N58), .E(N100), .CP(clk), .Q(\entry[7][8] ) );
  EDFQD1 \entry_reg[7][7]  ( .D(N57), .E(N100), .CP(clk), .Q(\entry[7][7] ) );
  EDFQD1 \entry_reg[7][6]  ( .D(N56), .E(N100), .CP(clk), .Q(\entry[7][6] ) );
  EDFQD1 \entry_reg[7][5]  ( .D(N55), .E(N100), .CP(clk), .Q(\entry[7][5] ) );
  EDFQD1 \entry_reg[7][4]  ( .D(N54), .E(N100), .CP(clk), .Q(\entry[7][4] ) );
  EDFQD1 \entry_reg[7][3]  ( .D(N53), .E(N100), .CP(clk), .Q(\entry[7][3] ) );
  EDFQD1 \entry_reg[7][2]  ( .D(N52), .E(N100), .CP(clk), .Q(\entry[7][2] ) );
  EDFQD1 \entry_reg[7][1]  ( .D(N51), .E(N100), .CP(clk), .Q(\entry[7][1] ) );
  EDFQD1 \entry_reg[7][0]  ( .D(N50), .E(N100), .CP(clk), .Q(\entry[7][0] ) );
  EDFQD1 \entry_reg[6][43]  ( .D(N93), .E(N99), .CP(clk), .Q(\entry[6][43] )
         );
  EDFQD1 \entry_reg[6][42]  ( .D(N92), .E(N99), .CP(clk), .Q(\entry[6][42] )
         );
  EDFQD1 \entry_reg[6][41]  ( .D(N91), .E(N99), .CP(clk), .Q(\entry[6][41] )
         );
  EDFQD1 \entry_reg[6][40]  ( .D(N90), .E(N99), .CP(clk), .Q(\entry[6][40] )
         );
  EDFQD1 \entry_reg[6][39]  ( .D(N89), .E(N99), .CP(clk), .Q(\entry[6][39] )
         );
  EDFQD1 \entry_reg[6][38]  ( .D(N88), .E(N99), .CP(clk), .Q(\entry[6][38] )
         );
  EDFQD1 \entry_reg[6][37]  ( .D(N87), .E(N99), .CP(clk), .Q(\entry[6][37] )
         );
  EDFQD1 \entry_reg[6][36]  ( .D(N86), .E(N99), .CP(clk), .Q(\entry[6][36] )
         );
  EDFQD1 \entry_reg[6][35]  ( .D(N85), .E(N99), .CP(clk), .Q(\entry[6][35] )
         );
  EDFQD1 \entry_reg[6][34]  ( .D(N84), .E(N99), .CP(clk), .Q(\entry[6][34] )
         );
  EDFQD1 \entry_reg[6][33]  ( .D(N83), .E(N99), .CP(clk), .Q(\entry[6][33] )
         );
  EDFQD1 \entry_reg[6][32]  ( .D(N82), .E(N99), .CP(clk), .Q(\entry[6][32] )
         );
  EDFQD1 \entry_reg[6][31]  ( .D(N81), .E(N99), .CP(clk), .Q(\entry[6][31] )
         );
  EDFQD1 \entry_reg[6][30]  ( .D(N80), .E(N99), .CP(clk), .Q(\entry[6][30] )
         );
  EDFQD1 \entry_reg[6][29]  ( .D(N79), .E(N99), .CP(clk), .Q(\entry[6][29] )
         );
  EDFQD1 \entry_reg[6][28]  ( .D(N78), .E(N99), .CP(clk), .Q(\entry[6][28] )
         );
  EDFQD1 \entry_reg[6][27]  ( .D(N77), .E(N99), .CP(clk), .Q(\entry[6][27] )
         );
  EDFQD1 \entry_reg[6][26]  ( .D(N76), .E(N99), .CP(clk), .Q(\entry[6][26] )
         );
  EDFQD1 \entry_reg[6][25]  ( .D(N75), .E(N99), .CP(clk), .Q(\entry[6][25] )
         );
  EDFQD1 \entry_reg[6][24]  ( .D(N74), .E(N99), .CP(clk), .Q(\entry[6][24] )
         );
  EDFQD1 \entry_reg[6][23]  ( .D(N73), .E(N99), .CP(clk), .Q(\entry[6][23] )
         );
  EDFQD1 \entry_reg[6][22]  ( .D(N72), .E(N99), .CP(clk), .Q(\entry[6][22] )
         );
  EDFQD1 \entry_reg[6][21]  ( .D(N71), .E(N99), .CP(clk), .Q(\entry[6][21] )
         );
  EDFQD1 \entry_reg[6][20]  ( .D(N70), .E(N99), .CP(clk), .Q(\entry[6][20] )
         );
  EDFQD1 \entry_reg[6][19]  ( .D(N69), .E(N99), .CP(clk), .Q(\entry[6][19] )
         );
  EDFQD1 \entry_reg[6][18]  ( .D(N68), .E(N99), .CP(clk), .Q(\entry[6][18] )
         );
  EDFQD1 \entry_reg[6][17]  ( .D(N67), .E(N99), .CP(clk), .Q(\entry[6][17] )
         );
  EDFQD1 \entry_reg[6][16]  ( .D(N66), .E(N99), .CP(clk), .Q(\entry[6][16] )
         );
  EDFQD1 \entry_reg[6][15]  ( .D(N65), .E(N99), .CP(clk), .Q(\entry[6][15] )
         );
  EDFQD1 \entry_reg[6][14]  ( .D(N64), .E(N99), .CP(clk), .Q(\entry[6][14] )
         );
  EDFQD1 \entry_reg[6][13]  ( .D(N63), .E(N99), .CP(clk), .Q(\entry[6][13] )
         );
  EDFQD1 \entry_reg[6][12]  ( .D(N62), .E(N99), .CP(clk), .Q(\entry[6][12] )
         );
  EDFQD1 \entry_reg[6][11]  ( .D(N61), .E(N99), .CP(clk), .Q(\entry[6][11] )
         );
  EDFQD1 \entry_reg[6][10]  ( .D(N60), .E(N99), .CP(clk), .Q(\entry[6][10] )
         );
  EDFQD1 \entry_reg[6][9]  ( .D(N59), .E(N99), .CP(clk), .Q(\entry[6][9] ) );
  EDFQD1 \entry_reg[6][8]  ( .D(N58), .E(N99), .CP(clk), .Q(\entry[6][8] ) );
  EDFQD1 \entry_reg[6][7]  ( .D(N57), .E(N99), .CP(clk), .Q(\entry[6][7] ) );
  EDFQD1 \entry_reg[6][6]  ( .D(N56), .E(N99), .CP(clk), .Q(\entry[6][6] ) );
  EDFQD1 \entry_reg[6][5]  ( .D(N55), .E(N99), .CP(clk), .Q(\entry[6][5] ) );
  EDFQD1 \entry_reg[6][4]  ( .D(N54), .E(N99), .CP(clk), .Q(\entry[6][4] ) );
  EDFQD1 \entry_reg[6][3]  ( .D(N53), .E(N99), .CP(clk), .Q(\entry[6][3] ) );
  EDFQD1 \entry_reg[6][2]  ( .D(N52), .E(N99), .CP(clk), .Q(\entry[6][2] ) );
  EDFQD1 \entry_reg[6][1]  ( .D(N51), .E(N99), .CP(clk), .Q(\entry[6][1] ) );
  EDFQD1 \entry_reg[6][0]  ( .D(N50), .E(N99), .CP(clk), .Q(\entry[6][0] ) );
  EDFQD1 \entry_reg[5][43]  ( .D(N93), .E(N98), .CP(clk), .Q(\entry[5][43] )
         );
  EDFQD1 \entry_reg[5][42]  ( .D(N92), .E(N98), .CP(clk), .Q(\entry[5][42] )
         );
  EDFQD1 \entry_reg[5][41]  ( .D(N91), .E(N98), .CP(clk), .Q(\entry[5][41] )
         );
  EDFQD1 \entry_reg[5][40]  ( .D(N90), .E(N98), .CP(clk), .Q(\entry[5][40] )
         );
  EDFQD1 \entry_reg[5][39]  ( .D(N89), .E(N98), .CP(clk), .Q(\entry[5][39] )
         );
  EDFQD1 \entry_reg[5][38]  ( .D(N88), .E(N98), .CP(clk), .Q(\entry[5][38] )
         );
  EDFQD1 \entry_reg[5][37]  ( .D(N87), .E(N98), .CP(clk), .Q(\entry[5][37] )
         );
  EDFQD1 \entry_reg[5][36]  ( .D(N86), .E(N98), .CP(clk), .Q(\entry[5][36] )
         );
  EDFQD1 \entry_reg[5][35]  ( .D(N85), .E(N98), .CP(clk), .Q(\entry[5][35] )
         );
  EDFQD1 \entry_reg[5][34]  ( .D(N84), .E(N98), .CP(clk), .Q(\entry[5][34] )
         );
  EDFQD1 \entry_reg[5][33]  ( .D(N83), .E(N98), .CP(clk), .Q(\entry[5][33] )
         );
  EDFQD1 \entry_reg[5][32]  ( .D(N82), .E(N98), .CP(clk), .Q(\entry[5][32] )
         );
  EDFQD1 \entry_reg[5][31]  ( .D(N81), .E(N98), .CP(clk), .Q(\entry[5][31] )
         );
  EDFQD1 \entry_reg[5][30]  ( .D(N80), .E(N98), .CP(clk), .Q(\entry[5][30] )
         );
  EDFQD1 \entry_reg[5][29]  ( .D(N79), .E(N98), .CP(clk), .Q(\entry[5][29] )
         );
  EDFQD1 \entry_reg[5][28]  ( .D(N78), .E(N98), .CP(clk), .Q(\entry[5][28] )
         );
  EDFQD1 \entry_reg[5][27]  ( .D(N77), .E(N98), .CP(clk), .Q(\entry[5][27] )
         );
  EDFQD1 \entry_reg[5][26]  ( .D(N76), .E(N98), .CP(clk), .Q(\entry[5][26] )
         );
  EDFQD1 \entry_reg[5][25]  ( .D(N75), .E(N98), .CP(clk), .Q(\entry[5][25] )
         );
  EDFQD1 \entry_reg[5][24]  ( .D(N74), .E(N98), .CP(clk), .Q(\entry[5][24] )
         );
  EDFQD1 \entry_reg[5][23]  ( .D(N73), .E(N98), .CP(clk), .Q(\entry[5][23] )
         );
  EDFQD1 \entry_reg[5][22]  ( .D(N72), .E(N98), .CP(clk), .Q(\entry[5][22] )
         );
  EDFQD1 \entry_reg[5][21]  ( .D(N71), .E(N98), .CP(clk), .Q(\entry[5][21] )
         );
  EDFQD1 \entry_reg[5][20]  ( .D(N70), .E(N98), .CP(clk), .Q(\entry[5][20] )
         );
  EDFQD1 \entry_reg[5][19]  ( .D(N69), .E(N98), .CP(clk), .Q(\entry[5][19] )
         );
  EDFQD1 \entry_reg[5][18]  ( .D(N68), .E(N98), .CP(clk), .Q(\entry[5][18] )
         );
  EDFQD1 \entry_reg[5][17]  ( .D(N67), .E(N98), .CP(clk), .Q(\entry[5][17] )
         );
  EDFQD1 \entry_reg[5][16]  ( .D(N66), .E(N98), .CP(clk), .Q(\entry[5][16] )
         );
  EDFQD1 \entry_reg[5][15]  ( .D(N65), .E(N98), .CP(clk), .Q(\entry[5][15] )
         );
  EDFQD1 \entry_reg[5][14]  ( .D(N64), .E(N98), .CP(clk), .Q(\entry[5][14] )
         );
  EDFQD1 \entry_reg[5][13]  ( .D(N63), .E(N98), .CP(clk), .Q(\entry[5][13] )
         );
  EDFQD1 \entry_reg[5][12]  ( .D(N62), .E(N98), .CP(clk), .Q(\entry[5][12] )
         );
  EDFQD1 \entry_reg[5][11]  ( .D(N61), .E(N98), .CP(clk), .Q(\entry[5][11] )
         );
  EDFQD1 \entry_reg[5][10]  ( .D(N60), .E(N98), .CP(clk), .Q(\entry[5][10] )
         );
  EDFQD1 \entry_reg[5][9]  ( .D(N59), .E(N98), .CP(clk), .Q(\entry[5][9] ) );
  EDFQD1 \entry_reg[5][8]  ( .D(N58), .E(N98), .CP(clk), .Q(\entry[5][8] ) );
  EDFQD1 \entry_reg[5][7]  ( .D(N57), .E(N98), .CP(clk), .Q(\entry[5][7] ) );
  EDFQD1 \entry_reg[5][6]  ( .D(N56), .E(N98), .CP(clk), .Q(\entry[5][6] ) );
  EDFQD1 \entry_reg[5][5]  ( .D(N55), .E(N98), .CP(clk), .Q(\entry[5][5] ) );
  EDFQD1 \entry_reg[5][4]  ( .D(N54), .E(N98), .CP(clk), .Q(\entry[5][4] ) );
  EDFQD1 \entry_reg[5][3]  ( .D(N53), .E(N98), .CP(clk), .Q(\entry[5][3] ) );
  EDFQD1 \entry_reg[5][2]  ( .D(N52), .E(N98), .CP(clk), .Q(\entry[5][2] ) );
  EDFQD1 \entry_reg[5][1]  ( .D(N51), .E(N98), .CP(clk), .Q(\entry[5][1] ) );
  EDFQD1 \entry_reg[5][0]  ( .D(N50), .E(N98), .CP(clk), .Q(\entry[5][0] ) );
  EDFQD1 \entry_reg[4][43]  ( .D(N93), .E(N97), .CP(clk), .Q(\entry[4][43] )
         );
  EDFQD1 \entry_reg[4][42]  ( .D(N92), .E(N97), .CP(clk), .Q(\entry[4][42] )
         );
  EDFQD1 \entry_reg[4][41]  ( .D(N91), .E(N97), .CP(clk), .Q(\entry[4][41] )
         );
  EDFQD1 \entry_reg[4][40]  ( .D(N90), .E(N97), .CP(clk), .Q(\entry[4][40] )
         );
  EDFQD1 \entry_reg[4][39]  ( .D(N89), .E(N97), .CP(clk), .Q(\entry[4][39] )
         );
  EDFQD1 \entry_reg[4][38]  ( .D(N88), .E(N97), .CP(clk), .Q(\entry[4][38] )
         );
  EDFQD1 \entry_reg[4][37]  ( .D(N87), .E(N97), .CP(clk), .Q(\entry[4][37] )
         );
  EDFQD1 \entry_reg[4][36]  ( .D(N86), .E(N97), .CP(clk), .Q(\entry[4][36] )
         );
  EDFQD1 \entry_reg[4][35]  ( .D(N85), .E(N97), .CP(clk), .Q(\entry[4][35] )
         );
  EDFQD1 \entry_reg[4][34]  ( .D(N84), .E(N97), .CP(clk), .Q(\entry[4][34] )
         );
  EDFQD1 \entry_reg[4][33]  ( .D(N83), .E(N97), .CP(clk), .Q(\entry[4][33] )
         );
  EDFQD1 \entry_reg[4][32]  ( .D(N82), .E(N97), .CP(clk), .Q(\entry[4][32] )
         );
  EDFQD1 \entry_reg[4][31]  ( .D(N81), .E(N97), .CP(clk), .Q(\entry[4][31] )
         );
  EDFQD1 \entry_reg[4][30]  ( .D(N80), .E(N97), .CP(clk), .Q(\entry[4][30] )
         );
  EDFQD1 \entry_reg[4][29]  ( .D(N79), .E(N97), .CP(clk), .Q(\entry[4][29] )
         );
  EDFQD1 \entry_reg[4][28]  ( .D(N78), .E(N97), .CP(clk), .Q(\entry[4][28] )
         );
  EDFQD1 \entry_reg[4][27]  ( .D(N77), .E(N97), .CP(clk), .Q(\entry[4][27] )
         );
  EDFQD1 \entry_reg[4][26]  ( .D(N76), .E(N97), .CP(clk), .Q(\entry[4][26] )
         );
  EDFQD1 \entry_reg[4][25]  ( .D(N75), .E(N97), .CP(clk), .Q(\entry[4][25] )
         );
  EDFQD1 \entry_reg[4][24]  ( .D(N74), .E(N97), .CP(clk), .Q(\entry[4][24] )
         );
  EDFQD1 \entry_reg[4][23]  ( .D(N73), .E(N97), .CP(clk), .Q(\entry[4][23] )
         );
  EDFQD1 \entry_reg[4][22]  ( .D(N72), .E(N97), .CP(clk), .Q(\entry[4][22] )
         );
  EDFQD1 \entry_reg[4][21]  ( .D(N71), .E(N97), .CP(clk), .Q(\entry[4][21] )
         );
  EDFQD1 \entry_reg[4][20]  ( .D(N70), .E(N97), .CP(clk), .Q(\entry[4][20] )
         );
  EDFQD1 \entry_reg[4][19]  ( .D(N69), .E(N97), .CP(clk), .Q(\entry[4][19] )
         );
  EDFQD1 \entry_reg[4][18]  ( .D(N68), .E(N97), .CP(clk), .Q(\entry[4][18] )
         );
  EDFQD1 \entry_reg[4][17]  ( .D(N67), .E(N97), .CP(clk), .Q(\entry[4][17] )
         );
  EDFQD1 \entry_reg[4][16]  ( .D(N66), .E(N97), .CP(clk), .Q(\entry[4][16] )
         );
  EDFQD1 \entry_reg[4][15]  ( .D(N65), .E(N97), .CP(clk), .Q(\entry[4][15] )
         );
  EDFQD1 \entry_reg[4][14]  ( .D(N64), .E(N97), .CP(clk), .Q(\entry[4][14] )
         );
  EDFQD1 \entry_reg[4][13]  ( .D(N63), .E(N97), .CP(clk), .Q(\entry[4][13] )
         );
  EDFQD1 \entry_reg[4][12]  ( .D(N62), .E(N97), .CP(clk), .Q(\entry[4][12] )
         );
  EDFQD1 \entry_reg[4][11]  ( .D(N61), .E(N97), .CP(clk), .Q(\entry[4][11] )
         );
  EDFQD1 \entry_reg[4][10]  ( .D(N60), .E(N97), .CP(clk), .Q(\entry[4][10] )
         );
  EDFQD1 \entry_reg[4][9]  ( .D(N59), .E(N97), .CP(clk), .Q(\entry[4][9] ) );
  EDFQD1 \entry_reg[4][8]  ( .D(N58), .E(N97), .CP(clk), .Q(\entry[4][8] ) );
  EDFQD1 \entry_reg[4][7]  ( .D(N57), .E(N97), .CP(clk), .Q(\entry[4][7] ) );
  EDFQD1 \entry_reg[4][6]  ( .D(N56), .E(N97), .CP(clk), .Q(\entry[4][6] ) );
  EDFQD1 \entry_reg[4][5]  ( .D(N55), .E(N97), .CP(clk), .Q(\entry[4][5] ) );
  EDFQD1 \entry_reg[4][4]  ( .D(N54), .E(N97), .CP(clk), .Q(\entry[4][4] ) );
  EDFQD1 \entry_reg[4][3]  ( .D(N53), .E(N97), .CP(clk), .Q(\entry[4][3] ) );
  EDFQD1 \entry_reg[4][2]  ( .D(N52), .E(N97), .CP(clk), .Q(\entry[4][2] ) );
  EDFQD1 \entry_reg[4][1]  ( .D(N51), .E(N97), .CP(clk), .Q(\entry[4][1] ) );
  EDFQD1 \entry_reg[4][0]  ( .D(N50), .E(N97), .CP(clk), .Q(\entry[4][0] ) );
  EDFQD1 \entry_reg[3][43]  ( .D(N93), .E(N96), .CP(clk), .Q(\entry[3][43] )
         );
  EDFQD1 \entry_reg[3][42]  ( .D(N92), .E(N96), .CP(clk), .Q(\entry[3][42] )
         );
  EDFQD1 \entry_reg[3][41]  ( .D(N91), .E(N96), .CP(clk), .Q(\entry[3][41] )
         );
  EDFQD1 \entry_reg[3][40]  ( .D(N90), .E(N96), .CP(clk), .Q(\entry[3][40] )
         );
  EDFQD1 \entry_reg[3][39]  ( .D(N89), .E(N96), .CP(clk), .Q(\entry[3][39] )
         );
  EDFQD1 \entry_reg[3][38]  ( .D(N88), .E(N96), .CP(clk), .Q(\entry[3][38] )
         );
  EDFQD1 \entry_reg[3][37]  ( .D(N87), .E(N96), .CP(clk), .Q(\entry[3][37] )
         );
  EDFQD1 \entry_reg[3][36]  ( .D(N86), .E(N96), .CP(clk), .Q(\entry[3][36] )
         );
  EDFQD1 \entry_reg[3][35]  ( .D(N85), .E(N96), .CP(clk), .Q(\entry[3][35] )
         );
  EDFQD1 \entry_reg[3][34]  ( .D(N84), .E(N96), .CP(clk), .Q(\entry[3][34] )
         );
  EDFQD1 \entry_reg[3][33]  ( .D(N83), .E(N96), .CP(clk), .Q(\entry[3][33] )
         );
  EDFQD1 \entry_reg[3][32]  ( .D(N82), .E(N96), .CP(clk), .Q(\entry[3][32] )
         );
  EDFQD1 \entry_reg[3][31]  ( .D(N81), .E(N96), .CP(clk), .Q(\entry[3][31] )
         );
  EDFQD1 \entry_reg[3][30]  ( .D(N80), .E(N96), .CP(clk), .Q(\entry[3][30] )
         );
  EDFQD1 \entry_reg[3][29]  ( .D(N79), .E(N96), .CP(clk), .Q(\entry[3][29] )
         );
  EDFQD1 \entry_reg[3][28]  ( .D(N78), .E(N96), .CP(clk), .Q(\entry[3][28] )
         );
  EDFQD1 \entry_reg[3][27]  ( .D(N77), .E(N96), .CP(clk), .Q(\entry[3][27] )
         );
  EDFQD1 \entry_reg[3][26]  ( .D(N76), .E(N96), .CP(clk), .Q(\entry[3][26] )
         );
  EDFQD1 \entry_reg[3][25]  ( .D(N75), .E(N96), .CP(clk), .Q(\entry[3][25] )
         );
  EDFQD1 \entry_reg[3][24]  ( .D(N74), .E(N96), .CP(clk), .Q(\entry[3][24] )
         );
  EDFQD1 \entry_reg[3][23]  ( .D(N73), .E(N96), .CP(clk), .Q(\entry[3][23] )
         );
  EDFQD1 \entry_reg[3][22]  ( .D(N72), .E(N96), .CP(clk), .Q(\entry[3][22] )
         );
  EDFQD1 \entry_reg[3][21]  ( .D(N71), .E(N96), .CP(clk), .Q(\entry[3][21] )
         );
  EDFQD1 \entry_reg[3][20]  ( .D(N70), .E(N96), .CP(clk), .Q(\entry[3][20] )
         );
  EDFQD1 \entry_reg[3][19]  ( .D(N69), .E(N96), .CP(clk), .Q(\entry[3][19] )
         );
  EDFQD1 \entry_reg[3][18]  ( .D(N68), .E(N96), .CP(clk), .Q(\entry[3][18] )
         );
  EDFQD1 \entry_reg[3][17]  ( .D(N67), .E(N96), .CP(clk), .Q(\entry[3][17] )
         );
  EDFQD1 \entry_reg[3][16]  ( .D(N66), .E(N96), .CP(clk), .Q(\entry[3][16] )
         );
  EDFQD1 \entry_reg[3][15]  ( .D(N65), .E(N96), .CP(clk), .Q(\entry[3][15] )
         );
  EDFQD1 \entry_reg[3][14]  ( .D(N64), .E(N96), .CP(clk), .Q(\entry[3][14] )
         );
  EDFQD1 \entry_reg[3][13]  ( .D(N63), .E(N96), .CP(clk), .Q(\entry[3][13] )
         );
  EDFQD1 \entry_reg[3][12]  ( .D(N62), .E(N96), .CP(clk), .Q(\entry[3][12] )
         );
  EDFQD1 \entry_reg[3][11]  ( .D(N61), .E(N96), .CP(clk), .Q(\entry[3][11] )
         );
  EDFQD1 \entry_reg[3][10]  ( .D(N60), .E(N96), .CP(clk), .Q(\entry[3][10] )
         );
  EDFQD1 \entry_reg[3][9]  ( .D(N59), .E(N96), .CP(clk), .Q(\entry[3][9] ) );
  EDFQD1 \entry_reg[3][8]  ( .D(N58), .E(N96), .CP(clk), .Q(\entry[3][8] ) );
  EDFQD1 \entry_reg[3][7]  ( .D(N57), .E(N96), .CP(clk), .Q(\entry[3][7] ) );
  EDFQD1 \entry_reg[3][6]  ( .D(N56), .E(N96), .CP(clk), .Q(\entry[3][6] ) );
  EDFQD1 \entry_reg[3][5]  ( .D(N55), .E(N96), .CP(clk), .Q(\entry[3][5] ) );
  EDFQD1 \entry_reg[3][4]  ( .D(N54), .E(N96), .CP(clk), .Q(\entry[3][4] ) );
  EDFQD1 \entry_reg[3][3]  ( .D(N53), .E(N96), .CP(clk), .Q(\entry[3][3] ) );
  EDFQD1 \entry_reg[3][2]  ( .D(N52), .E(N96), .CP(clk), .Q(\entry[3][2] ) );
  EDFQD1 \entry_reg[3][1]  ( .D(N51), .E(N96), .CP(clk), .Q(\entry[3][1] ) );
  EDFQD1 \entry_reg[3][0]  ( .D(N50), .E(N96), .CP(clk), .Q(\entry[3][0] ) );
  EDFQD1 \entry_reg[2][43]  ( .D(N93), .E(N95), .CP(clk), .Q(\entry[2][43] )
         );
  EDFQD1 \entry_reg[2][42]  ( .D(N92), .E(N95), .CP(clk), .Q(\entry[2][42] )
         );
  EDFQD1 \entry_reg[2][41]  ( .D(N91), .E(N95), .CP(clk), .Q(\entry[2][41] )
         );
  EDFQD1 \entry_reg[2][40]  ( .D(N90), .E(N95), .CP(clk), .Q(\entry[2][40] )
         );
  EDFQD1 \entry_reg[2][39]  ( .D(N89), .E(N95), .CP(clk), .Q(\entry[2][39] )
         );
  EDFQD1 \entry_reg[2][38]  ( .D(N88), .E(N95), .CP(clk), .Q(\entry[2][38] )
         );
  EDFQD1 \entry_reg[2][37]  ( .D(N87), .E(N95), .CP(clk), .Q(\entry[2][37] )
         );
  EDFQD1 \entry_reg[2][36]  ( .D(N86), .E(N95), .CP(clk), .Q(\entry[2][36] )
         );
  EDFQD1 \entry_reg[2][35]  ( .D(N85), .E(N95), .CP(clk), .Q(\entry[2][35] )
         );
  EDFQD1 \entry_reg[2][34]  ( .D(N84), .E(N95), .CP(clk), .Q(\entry[2][34] )
         );
  EDFQD1 \entry_reg[2][33]  ( .D(N83), .E(N95), .CP(clk), .Q(\entry[2][33] )
         );
  EDFQD1 \entry_reg[2][32]  ( .D(N82), .E(N95), .CP(clk), .Q(\entry[2][32] )
         );
  EDFQD1 \entry_reg[2][31]  ( .D(N81), .E(N95), .CP(clk), .Q(\entry[2][31] )
         );
  EDFQD1 \entry_reg[2][30]  ( .D(N80), .E(N95), .CP(clk), .Q(\entry[2][30] )
         );
  EDFQD1 \entry_reg[2][29]  ( .D(N79), .E(N95), .CP(clk), .Q(\entry[2][29] )
         );
  EDFQD1 \entry_reg[2][28]  ( .D(N78), .E(N95), .CP(clk), .Q(\entry[2][28] )
         );
  EDFQD1 \entry_reg[2][27]  ( .D(N77), .E(N95), .CP(clk), .Q(\entry[2][27] )
         );
  EDFQD1 \entry_reg[2][26]  ( .D(N76), .E(N95), .CP(clk), .Q(\entry[2][26] )
         );
  EDFQD1 \entry_reg[2][25]  ( .D(N75), .E(N95), .CP(clk), .Q(\entry[2][25] )
         );
  EDFQD1 \entry_reg[2][24]  ( .D(N74), .E(N95), .CP(clk), .Q(\entry[2][24] )
         );
  EDFQD1 \entry_reg[2][23]  ( .D(N73), .E(N95), .CP(clk), .Q(\entry[2][23] )
         );
  EDFQD1 \entry_reg[2][22]  ( .D(N72), .E(N95), .CP(clk), .Q(\entry[2][22] )
         );
  EDFQD1 \entry_reg[2][21]  ( .D(N71), .E(N95), .CP(clk), .Q(\entry[2][21] )
         );
  EDFQD1 \entry_reg[2][20]  ( .D(N70), .E(N95), .CP(clk), .Q(\entry[2][20] )
         );
  EDFQD1 \entry_reg[2][19]  ( .D(N69), .E(N95), .CP(clk), .Q(\entry[2][19] )
         );
  EDFQD1 \entry_reg[2][18]  ( .D(N68), .E(N95), .CP(clk), .Q(\entry[2][18] )
         );
  EDFQD1 \entry_reg[2][17]  ( .D(N67), .E(N95), .CP(clk), .Q(\entry[2][17] )
         );
  EDFQD1 \entry_reg[2][16]  ( .D(N66), .E(N95), .CP(clk), .Q(\entry[2][16] )
         );
  EDFQD1 \entry_reg[2][15]  ( .D(N65), .E(N95), .CP(clk), .Q(\entry[2][15] )
         );
  EDFQD1 \entry_reg[2][14]  ( .D(N64), .E(N95), .CP(clk), .Q(\entry[2][14] )
         );
  EDFQD1 \entry_reg[2][13]  ( .D(N63), .E(N95), .CP(clk), .Q(\entry[2][13] )
         );
  EDFQD1 \entry_reg[2][12]  ( .D(N62), .E(N95), .CP(clk), .Q(\entry[2][12] )
         );
  EDFQD1 \entry_reg[2][11]  ( .D(N61), .E(N95), .CP(clk), .Q(\entry[2][11] )
         );
  EDFQD1 \entry_reg[2][10]  ( .D(N60), .E(N95), .CP(clk), .Q(\entry[2][10] )
         );
  EDFQD1 \entry_reg[2][9]  ( .D(N59), .E(N95), .CP(clk), .Q(\entry[2][9] ) );
  EDFQD1 \entry_reg[2][8]  ( .D(N58), .E(N95), .CP(clk), .Q(\entry[2][8] ) );
  EDFQD1 \entry_reg[2][7]  ( .D(N57), .E(N95), .CP(clk), .Q(\entry[2][7] ) );
  EDFQD1 \entry_reg[2][6]  ( .D(N56), .E(N95), .CP(clk), .Q(\entry[2][6] ) );
  EDFQD1 \entry_reg[2][5]  ( .D(N55), .E(N95), .CP(clk), .Q(\entry[2][5] ) );
  EDFQD1 \entry_reg[2][4]  ( .D(N54), .E(N95), .CP(clk), .Q(\entry[2][4] ) );
  EDFQD1 \entry_reg[2][3]  ( .D(N53), .E(N95), .CP(clk), .Q(\entry[2][3] ) );
  EDFQD1 \entry_reg[2][2]  ( .D(N52), .E(N95), .CP(clk), .Q(\entry[2][2] ) );
  EDFQD1 \entry_reg[2][1]  ( .D(N51), .E(N95), .CP(clk), .Q(\entry[2][1] ) );
  EDFQD1 \entry_reg[2][0]  ( .D(N50), .E(N95), .CP(clk), .Q(\entry[2][0] ) );
  EDFQD1 \entry_reg[1][43]  ( .D(N93), .E(N94), .CP(clk), .Q(\entry[1][43] )
         );
  EDFQD1 \entry_reg[1][42]  ( .D(N92), .E(N94), .CP(clk), .Q(\entry[1][42] )
         );
  EDFQD1 \entry_reg[1][41]  ( .D(N91), .E(N94), .CP(clk), .Q(\entry[1][41] )
         );
  EDFQD1 \entry_reg[1][40]  ( .D(N90), .E(N94), .CP(clk), .Q(\entry[1][40] )
         );
  EDFQD1 \entry_reg[1][39]  ( .D(N89), .E(N94), .CP(clk), .Q(\entry[1][39] )
         );
  EDFQD1 \entry_reg[1][38]  ( .D(N88), .E(N94), .CP(clk), .Q(\entry[1][38] )
         );
  EDFQD1 \entry_reg[1][37]  ( .D(N87), .E(N94), .CP(clk), .Q(\entry[1][37] )
         );
  EDFQD1 \entry_reg[1][36]  ( .D(N86), .E(N94), .CP(clk), .Q(\entry[1][36] )
         );
  EDFQD1 \entry_reg[1][35]  ( .D(N85), .E(N94), .CP(clk), .Q(\entry[1][35] )
         );
  EDFQD1 \entry_reg[1][34]  ( .D(N84), .E(N94), .CP(clk), .Q(\entry[1][34] )
         );
  EDFQD1 \entry_reg[1][33]  ( .D(N83), .E(N94), .CP(clk), .Q(\entry[1][33] )
         );
  EDFQD1 \entry_reg[1][32]  ( .D(N82), .E(N94), .CP(clk), .Q(\entry[1][32] )
         );
  EDFQD1 \entry_reg[1][31]  ( .D(N81), .E(N94), .CP(clk), .Q(\entry[1][31] )
         );
  EDFQD1 \entry_reg[1][30]  ( .D(N80), .E(N94), .CP(clk), .Q(\entry[1][30] )
         );
  EDFQD1 \entry_reg[1][29]  ( .D(N79), .E(N94), .CP(clk), .Q(\entry[1][29] )
         );
  EDFQD1 \entry_reg[1][28]  ( .D(N78), .E(N94), .CP(clk), .Q(\entry[1][28] )
         );
  EDFQD1 \entry_reg[1][27]  ( .D(N77), .E(N94), .CP(clk), .Q(\entry[1][27] )
         );
  EDFQD1 \entry_reg[1][26]  ( .D(N76), .E(N94), .CP(clk), .Q(\entry[1][26] )
         );
  EDFQD1 \entry_reg[1][25]  ( .D(N75), .E(N94), .CP(clk), .Q(\entry[1][25] )
         );
  EDFQD1 \entry_reg[1][24]  ( .D(N74), .E(N94), .CP(clk), .Q(\entry[1][24] )
         );
  EDFQD1 \entry_reg[1][23]  ( .D(N73), .E(N94), .CP(clk), .Q(\entry[1][23] )
         );
  EDFQD1 \entry_reg[1][22]  ( .D(N72), .E(N94), .CP(clk), .Q(\entry[1][22] )
         );
  EDFQD1 \entry_reg[1][21]  ( .D(N71), .E(N94), .CP(clk), .Q(\entry[1][21] )
         );
  EDFQD1 \entry_reg[1][20]  ( .D(N70), .E(N94), .CP(clk), .Q(\entry[1][20] )
         );
  EDFQD1 \entry_reg[1][19]  ( .D(N69), .E(N94), .CP(clk), .Q(\entry[1][19] )
         );
  EDFQD1 \entry_reg[1][18]  ( .D(N68), .E(N94), .CP(clk), .Q(\entry[1][18] )
         );
  EDFQD1 \entry_reg[1][17]  ( .D(N67), .E(N94), .CP(clk), .Q(\entry[1][17] )
         );
  EDFQD1 \entry_reg[1][16]  ( .D(N66), .E(N94), .CP(clk), .Q(\entry[1][16] )
         );
  EDFQD1 \entry_reg[1][15]  ( .D(N65), .E(N94), .CP(clk), .Q(\entry[1][15] )
         );
  EDFQD1 \entry_reg[1][14]  ( .D(N64), .E(N94), .CP(clk), .Q(\entry[1][14] )
         );
  EDFQD1 \entry_reg[1][13]  ( .D(N63), .E(N94), .CP(clk), .Q(\entry[1][13] )
         );
  EDFQD1 \entry_reg[1][12]  ( .D(N62), .E(N94), .CP(clk), .Q(\entry[1][12] )
         );
  EDFQD1 \entry_reg[1][11]  ( .D(N61), .E(N94), .CP(clk), .Q(\entry[1][11] )
         );
  EDFQD1 \entry_reg[1][10]  ( .D(N60), .E(N94), .CP(clk), .Q(\entry[1][10] )
         );
  EDFQD1 \entry_reg[1][9]  ( .D(N59), .E(N94), .CP(clk), .Q(\entry[1][9] ) );
  EDFQD1 \entry_reg[1][8]  ( .D(N58), .E(N94), .CP(clk), .Q(\entry[1][8] ) );
  EDFQD1 \entry_reg[1][7]  ( .D(N57), .E(N94), .CP(clk), .Q(\entry[1][7] ) );
  EDFQD1 \entry_reg[1][6]  ( .D(N56), .E(N94), .CP(clk), .Q(\entry[1][6] ) );
  EDFQD1 \entry_reg[1][5]  ( .D(N55), .E(N94), .CP(clk), .Q(\entry[1][5] ) );
  EDFQD1 \entry_reg[1][4]  ( .D(N54), .E(N94), .CP(clk), .Q(\entry[1][4] ) );
  EDFQD1 \entry_reg[1][3]  ( .D(N53), .E(N94), .CP(clk), .Q(\entry[1][3] ) );
  EDFQD1 \entry_reg[1][2]  ( .D(N52), .E(N94), .CP(clk), .Q(\entry[1][2] ) );
  EDFQD1 \entry_reg[1][1]  ( .D(N51), .E(N94), .CP(clk), .Q(\entry[1][1] ) );
  EDFQD1 \entry_reg[1][0]  ( .D(N50), .E(N94), .CP(clk), .Q(\entry[1][0] ) );
  EDFQD1 \entry_reg[0][43]  ( .D(N93), .E(N49), .CP(clk), .Q(\entry[0][43] )
         );
  EDFQD1 \entry_reg[0][42]  ( .D(N92), .E(N49), .CP(clk), .Q(\entry[0][42] )
         );
  EDFQD1 \entry_reg[0][41]  ( .D(N91), .E(N49), .CP(clk), .Q(\entry[0][41] )
         );
  EDFQD1 \entry_reg[0][40]  ( .D(N90), .E(N49), .CP(clk), .Q(\entry[0][40] )
         );
  EDFQD1 \entry_reg[0][39]  ( .D(N89), .E(N49), .CP(clk), .Q(\entry[0][39] )
         );
  EDFQD1 \entry_reg[0][38]  ( .D(N88), .E(N49), .CP(clk), .Q(\entry[0][38] )
         );
  EDFQD1 \entry_reg[0][37]  ( .D(N87), .E(N49), .CP(clk), .Q(\entry[0][37] )
         );
  EDFQD1 \entry_reg[0][36]  ( .D(N86), .E(N49), .CP(clk), .Q(\entry[0][36] )
         );
  EDFQD1 \entry_reg[0][35]  ( .D(N85), .E(N49), .CP(clk), .Q(\entry[0][35] )
         );
  EDFQD1 \entry_reg[0][34]  ( .D(N84), .E(N49), .CP(clk), .Q(\entry[0][34] )
         );
  EDFQD1 \entry_reg[0][33]  ( .D(N83), .E(N49), .CP(clk), .Q(\entry[0][33] )
         );
  EDFQD1 \entry_reg[0][32]  ( .D(N82), .E(N49), .CP(clk), .Q(\entry[0][32] )
         );
  EDFQD1 \entry_reg[0][31]  ( .D(N81), .E(N49), .CP(clk), .Q(\entry[0][31] )
         );
  EDFQD1 \entry_reg[0][30]  ( .D(N80), .E(N49), .CP(clk), .Q(\entry[0][30] )
         );
  EDFQD1 \entry_reg[0][29]  ( .D(N79), .E(N49), .CP(clk), .Q(\entry[0][29] )
         );
  EDFQD1 \entry_reg[0][28]  ( .D(N78), .E(N49), .CP(clk), .Q(\entry[0][28] )
         );
  EDFQD1 \entry_reg[0][27]  ( .D(N77), .E(N49), .CP(clk), .Q(\entry[0][27] )
         );
  EDFQD1 \entry_reg[0][26]  ( .D(N76), .E(N49), .CP(clk), .Q(\entry[0][26] )
         );
  EDFQD1 \entry_reg[0][25]  ( .D(N75), .E(N49), .CP(clk), .Q(\entry[0][25] )
         );
  EDFQD1 \entry_reg[0][24]  ( .D(N74), .E(N49), .CP(clk), .Q(\entry[0][24] )
         );
  EDFQD1 \entry_reg[0][23]  ( .D(N73), .E(N49), .CP(clk), .Q(\entry[0][23] )
         );
  EDFQD1 \entry_reg[0][22]  ( .D(N72), .E(N49), .CP(clk), .Q(\entry[0][22] )
         );
  EDFQD1 \entry_reg[0][21]  ( .D(N71), .E(N49), .CP(clk), .Q(\entry[0][21] )
         );
  EDFQD1 \entry_reg[0][20]  ( .D(N70), .E(N49), .CP(clk), .Q(\entry[0][20] )
         );
  EDFQD1 \entry_reg[0][19]  ( .D(N69), .E(N49), .CP(clk), .Q(\entry[0][19] )
         );
  EDFQD1 \entry_reg[0][18]  ( .D(N68), .E(N49), .CP(clk), .Q(\entry[0][18] )
         );
  EDFQD1 \entry_reg[0][17]  ( .D(N67), .E(N49), .CP(clk), .Q(\entry[0][17] )
         );
  EDFQD1 \entry_reg[0][16]  ( .D(N66), .E(N49), .CP(clk), .Q(\entry[0][16] )
         );
  EDFQD1 \entry_reg[0][15]  ( .D(N65), .E(N49), .CP(clk), .Q(\entry[0][15] )
         );
  EDFQD1 \entry_reg[0][14]  ( .D(N64), .E(N49), .CP(clk), .Q(\entry[0][14] )
         );
  EDFQD1 \entry_reg[0][13]  ( .D(N63), .E(N49), .CP(clk), .Q(\entry[0][13] )
         );
  EDFQD1 \entry_reg[0][12]  ( .D(N62), .E(N49), .CP(clk), .Q(\entry[0][12] )
         );
  EDFQD1 \entry_reg[0][11]  ( .D(N61), .E(N49), .CP(clk), .Q(\entry[0][11] )
         );
  EDFQD1 \entry_reg[0][10]  ( .D(N60), .E(N49), .CP(clk), .Q(\entry[0][10] )
         );
  EDFQD1 \entry_reg[0][9]  ( .D(N59), .E(N49), .CP(clk), .Q(\entry[0][9] ) );
  EDFQD1 \entry_reg[0][8]  ( .D(N58), .E(N49), .CP(clk), .Q(\entry[0][8] ) );
  EDFQD1 \entry_reg[0][7]  ( .D(N57), .E(N49), .CP(clk), .Q(\entry[0][7] ) );
  EDFQD1 \entry_reg[0][6]  ( .D(N56), .E(N49), .CP(clk), .Q(\entry[0][6] ) );
  EDFQD1 \entry_reg[0][5]  ( .D(N55), .E(N49), .CP(clk), .Q(\entry[0][5] ) );
  EDFQD1 \entry_reg[0][4]  ( .D(N54), .E(N49), .CP(clk), .Q(\entry[0][4] ) );
  EDFQD1 \entry_reg[0][3]  ( .D(N53), .E(N49), .CP(clk), .Q(\entry[0][3] ) );
  EDFQD1 \entry_reg[0][2]  ( .D(N52), .E(N49), .CP(clk), .Q(\entry[0][2] ) );
  EDFQD1 \entry_reg[0][1]  ( .D(N51), .E(N49), .CP(clk), .Q(\entry[0][1] ) );
  EDFQD1 \entry_reg[0][0]  ( .D(N50), .E(N49), .CP(clk), .Q(\entry[0][0] ) );
  ND2D1 U545 ( .A1(n587), .A2(n590), .ZN(N96) );
  OR2D1 U546 ( .A1(n779), .A2(count[2]), .Z(n590) );
  OAI21D2 U547 ( .A1(n588), .A2(n589), .B(n587), .ZN(N98) );
  OAI21D2 U548 ( .A1(count[2]), .A2(n589), .B(n587), .ZN(N94) );
  OAI21D2 U549 ( .A1(n585), .A2(n586), .B(n587), .ZN(N99) );
  OAI21D2 U550 ( .A1(n588), .A2(n779), .B(n587), .ZN(N100) );
  OAI21D2 U551 ( .A1(count[1]), .A2(n585), .B(n587), .ZN(N97) );
  OAI31D4 U552 ( .A1(n586), .A2(count[2]), .A3(n591), .B(n587), .ZN(N95) );
  ND4D1 U553 ( .A1(n682), .A2(n681), .A3(n683), .A4(n684), .ZN(N105) );
  OAI31D4 U554 ( .A1(n591), .A2(count[2]), .A3(count[1]), .B(n587), .ZN(N49)
         );
  INR2D0 U555 ( .A1(tag[23]), .B1(n592), .ZN(N93) );
  INR2D0 U556 ( .A1(tag[22]), .B1(n592), .ZN(N92) );
  INR2D0 U557 ( .A1(tag[21]), .B1(n592), .ZN(N91) );
  INR2D0 U558 ( .A1(tag[20]), .B1(n592), .ZN(N90) );
  INR2D0 U559 ( .A1(tag[19]), .B1(n592), .ZN(N89) );
  INR2D0 U560 ( .A1(tag[18]), .B1(n592), .ZN(N88) );
  INR2D0 U561 ( .A1(tag[17]), .B1(n592), .ZN(N87) );
  INR2D0 U562 ( .A1(tag[16]), .B1(n592), .ZN(N86) );
  INR2D0 U563 ( .A1(tag[15]), .B1(n592), .ZN(N85) );
  INR2D0 U564 ( .A1(tag[14]), .B1(n592), .ZN(N84) );
  INR2D0 U565 ( .A1(tag[13]), .B1(n592), .ZN(N83) );
  INR2D0 U566 ( .A1(tag[12]), .B1(n592), .ZN(N82) );
  INR2D0 U567 ( .A1(tag[11]), .B1(n592), .ZN(N81) );
  INR2D0 U568 ( .A1(tag[10]), .B1(n592), .ZN(N80) );
  INR2D0 U569 ( .A1(tag[9]), .B1(n592), .ZN(N79) );
  INR2D0 U570 ( .A1(tag[8]), .B1(n592), .ZN(N78) );
  INR2D0 U571 ( .A1(tag[7]), .B1(n592), .ZN(N77) );
  INR2D0 U572 ( .A1(tag[6]), .B1(n592), .ZN(N76) );
  INR2D0 U573 ( .A1(tag[5]), .B1(n592), .ZN(N75) );
  INR2D0 U574 ( .A1(tag[4]), .B1(n592), .ZN(N74) );
  INR2D0 U575 ( .A1(tag[3]), .B1(n592), .ZN(N73) );
  INR2D0 U576 ( .A1(tag[2]), .B1(n592), .ZN(N72) );
  INR2D0 U577 ( .A1(tag[1]), .B1(n592), .ZN(N71) );
  INR2D0 U578 ( .A1(tag[0]), .B1(n592), .ZN(N70) );
  INR2D0 U579 ( .A1(val[19]), .B1(n592), .ZN(N69) );
  INR2D0 U580 ( .A1(val[18]), .B1(n592), .ZN(N68) );
  INR2D0 U581 ( .A1(val[17]), .B1(n592), .ZN(N67) );
  INR2D0 U582 ( .A1(val[16]), .B1(n592), .ZN(N66) );
  INR2D0 U583 ( .A1(val[15]), .B1(n592), .ZN(N65) );
  INR2D0 U584 ( .A1(val[14]), .B1(n592), .ZN(N64) );
  INR2D0 U585 ( .A1(val[13]), .B1(n592), .ZN(N63) );
  INR2D0 U586 ( .A1(val[12]), .B1(n592), .ZN(N62) );
  INR2D0 U587 ( .A1(val[11]), .B1(n592), .ZN(N61) );
  INR2D0 U588 ( .A1(val[10]), .B1(n592), .ZN(N60) );
  INR2D0 U589 ( .A1(val[9]), .B1(n592), .ZN(N59) );
  INR2D0 U590 ( .A1(val[8]), .B1(n592), .ZN(N58) );
  INR2D0 U591 ( .A1(val[7]), .B1(n592), .ZN(N57) );
  INR2D0 U592 ( .A1(val[6]), .B1(n592), .ZN(N56) );
  INR2D0 U593 ( .A1(val[5]), .B1(n592), .ZN(N55) );
  INR2D0 U594 ( .A1(val[4]), .B1(n592), .ZN(N54) );
  INR2D0 U595 ( .A1(val[3]), .B1(n592), .ZN(N53) );
  INR2D0 U596 ( .A1(val[2]), .B1(n592), .ZN(N52) );
  INR2D0 U597 ( .A1(val[1]), .B1(n592), .ZN(N51) );
  INR2D0 U598 ( .A1(val[0]), .B1(n592), .ZN(N50) );
  ND4D0 U599 ( .A1(n593), .A2(n594), .A3(n595), .A4(n596), .ZN(N125) );
  AOI22D0 U600 ( .A1(\entry[2][19] ), .A2(n597), .B1(\entry[3][19] ), .B2(n598), .ZN(n596) );
  AOI22D0 U601 ( .A1(\entry[0][19] ), .A2(n599), .B1(\entry[5][19] ), .B2(n600), .ZN(n595) );
  AOI22D0 U602 ( .A1(\entry[1][19] ), .A2(n601), .B1(\entry[7][19] ), .B2(n602), .ZN(n594) );
  AOI22D0 U603 ( .A1(\entry[6][19] ), .A2(n603), .B1(\entry[4][19] ), .B2(n604), .ZN(n593) );
  ND4D0 U604 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(N124) );
  AOI22D0 U605 ( .A1(\entry[2][18] ), .A2(n597), .B1(\entry[3][18] ), .B2(n598), .ZN(n608) );
  AOI22D0 U606 ( .A1(\entry[0][18] ), .A2(n599), .B1(\entry[5][18] ), .B2(n600), .ZN(n607) );
  AOI22D0 U607 ( .A1(\entry[1][18] ), .A2(n601), .B1(\entry[7][18] ), .B2(n602), .ZN(n606) );
  AOI22D0 U608 ( .A1(\entry[6][18] ), .A2(n603), .B1(\entry[4][18] ), .B2(n604), .ZN(n605) );
  ND4D0 U609 ( .A1(n609), .A2(n610), .A3(n611), .A4(n612), .ZN(N123) );
  AOI22D0 U610 ( .A1(\entry[2][17] ), .A2(n597), .B1(\entry[3][17] ), .B2(n598), .ZN(n612) );
  AOI22D0 U611 ( .A1(\entry[0][17] ), .A2(n599), .B1(\entry[5][17] ), .B2(n600), .ZN(n611) );
  AOI22D0 U612 ( .A1(\entry[1][17] ), .A2(n601), .B1(\entry[7][17] ), .B2(n602), .ZN(n610) );
  AOI22D0 U613 ( .A1(\entry[6][17] ), .A2(n603), .B1(\entry[4][17] ), .B2(n604), .ZN(n609) );
  ND4D0 U614 ( .A1(n613), .A2(n614), .A3(n615), .A4(n616), .ZN(N122) );
  AOI22D0 U615 ( .A1(\entry[2][16] ), .A2(n597), .B1(\entry[3][16] ), .B2(n598), .ZN(n616) );
  AOI22D0 U616 ( .A1(\entry[0][16] ), .A2(n599), .B1(\entry[5][16] ), .B2(n600), .ZN(n615) );
  AOI22D0 U617 ( .A1(\entry[1][16] ), .A2(n601), .B1(\entry[7][16] ), .B2(n602), .ZN(n614) );
  AOI22D0 U618 ( .A1(\entry[6][16] ), .A2(n603), .B1(\entry[4][16] ), .B2(n604), .ZN(n613) );
  ND4D0 U619 ( .A1(n617), .A2(n618), .A3(n619), .A4(n620), .ZN(N121) );
  AOI22D0 U620 ( .A1(\entry[2][15] ), .A2(n597), .B1(\entry[3][15] ), .B2(n598), .ZN(n620) );
  AOI22D0 U621 ( .A1(\entry[0][15] ), .A2(n599), .B1(\entry[5][15] ), .B2(n600), .ZN(n619) );
  AOI22D0 U622 ( .A1(\entry[1][15] ), .A2(n601), .B1(\entry[7][15] ), .B2(n602), .ZN(n618) );
  AOI22D0 U623 ( .A1(\entry[6][15] ), .A2(n603), .B1(\entry[4][15] ), .B2(n604), .ZN(n617) );
  ND4D0 U624 ( .A1(n621), .A2(n622), .A3(n623), .A4(n624), .ZN(N120) );
  AOI22D0 U625 ( .A1(\entry[2][14] ), .A2(n597), .B1(\entry[3][14] ), .B2(n598), .ZN(n624) );
  AOI22D0 U626 ( .A1(\entry[0][14] ), .A2(n599), .B1(\entry[5][14] ), .B2(n600), .ZN(n623) );
  AOI22D0 U627 ( .A1(\entry[1][14] ), .A2(n601), .B1(\entry[7][14] ), .B2(n602), .ZN(n622) );
  AOI22D0 U628 ( .A1(\entry[6][14] ), .A2(n603), .B1(\entry[4][14] ), .B2(n604), .ZN(n621) );
  ND4D0 U629 ( .A1(n625), .A2(n626), .A3(n627), .A4(n628), .ZN(N119) );
  AOI22D0 U630 ( .A1(\entry[2][13] ), .A2(n597), .B1(\entry[3][13] ), .B2(n598), .ZN(n628) );
  AOI22D0 U631 ( .A1(\entry[0][13] ), .A2(n599), .B1(\entry[5][13] ), .B2(n600), .ZN(n627) );
  AOI22D0 U632 ( .A1(\entry[1][13] ), .A2(n601), .B1(\entry[7][13] ), .B2(n602), .ZN(n626) );
  AOI22D0 U633 ( .A1(\entry[6][13] ), .A2(n603), .B1(\entry[4][13] ), .B2(n604), .ZN(n625) );
  ND4D0 U634 ( .A1(n629), .A2(n630), .A3(n631), .A4(n632), .ZN(N118) );
  AOI22D0 U635 ( .A1(\entry[2][12] ), .A2(n597), .B1(\entry[3][12] ), .B2(n598), .ZN(n632) );
  AOI22D0 U636 ( .A1(\entry[0][12] ), .A2(n599), .B1(\entry[5][12] ), .B2(n600), .ZN(n631) );
  AOI22D0 U637 ( .A1(\entry[1][12] ), .A2(n601), .B1(\entry[7][12] ), .B2(n602), .ZN(n630) );
  AOI22D0 U638 ( .A1(\entry[6][12] ), .A2(n603), .B1(\entry[4][12] ), .B2(n604), .ZN(n629) );
  ND4D0 U639 ( .A1(n633), .A2(n634), .A3(n635), .A4(n636), .ZN(N117) );
  AOI22D0 U640 ( .A1(\entry[2][11] ), .A2(n597), .B1(\entry[3][11] ), .B2(n598), .ZN(n636) );
  AOI22D0 U641 ( .A1(\entry[0][11] ), .A2(n599), .B1(\entry[5][11] ), .B2(n600), .ZN(n635) );
  AOI22D0 U642 ( .A1(\entry[1][11] ), .A2(n601), .B1(\entry[7][11] ), .B2(n602), .ZN(n634) );
  AOI22D0 U643 ( .A1(\entry[6][11] ), .A2(n603), .B1(\entry[4][11] ), .B2(n604), .ZN(n633) );
  ND4D0 U644 ( .A1(n637), .A2(n638), .A3(n639), .A4(n640), .ZN(N116) );
  AOI22D0 U645 ( .A1(\entry[2][10] ), .A2(n597), .B1(\entry[3][10] ), .B2(n598), .ZN(n640) );
  AOI22D0 U646 ( .A1(\entry[0][10] ), .A2(n599), .B1(\entry[5][10] ), .B2(n600), .ZN(n639) );
  AOI22D0 U647 ( .A1(\entry[1][10] ), .A2(n601), .B1(\entry[7][10] ), .B2(n602), .ZN(n638) );
  AOI22D0 U648 ( .A1(\entry[6][10] ), .A2(n603), .B1(\entry[4][10] ), .B2(n604), .ZN(n637) );
  ND4D0 U649 ( .A1(n641), .A2(n642), .A3(n643), .A4(n644), .ZN(N115) );
  AOI22D0 U650 ( .A1(\entry[2][9] ), .A2(n597), .B1(\entry[3][9] ), .B2(n598), 
        .ZN(n644) );
  AOI22D0 U651 ( .A1(\entry[0][9] ), .A2(n599), .B1(\entry[5][9] ), .B2(n600), 
        .ZN(n643) );
  AOI22D0 U652 ( .A1(\entry[1][9] ), .A2(n601), .B1(\entry[7][9] ), .B2(n602), 
        .ZN(n642) );
  AOI22D0 U653 ( .A1(\entry[6][9] ), .A2(n603), .B1(\entry[4][9] ), .B2(n604), 
        .ZN(n641) );
  ND4D0 U654 ( .A1(n645), .A2(n646), .A3(n647), .A4(n648), .ZN(N114) );
  AOI22D0 U655 ( .A1(\entry[2][8] ), .A2(n597), .B1(\entry[3][8] ), .B2(n598), 
        .ZN(n648) );
  AOI22D0 U656 ( .A1(\entry[0][8] ), .A2(n599), .B1(\entry[5][8] ), .B2(n600), 
        .ZN(n647) );
  AOI22D0 U657 ( .A1(\entry[1][8] ), .A2(n601), .B1(\entry[7][8] ), .B2(n602), 
        .ZN(n646) );
  AOI22D0 U658 ( .A1(\entry[6][8] ), .A2(n603), .B1(\entry[4][8] ), .B2(n604), 
        .ZN(n645) );
  ND4D0 U659 ( .A1(n649), .A2(n650), .A3(n651), .A4(n652), .ZN(N113) );
  AOI22D0 U660 ( .A1(\entry[2][7] ), .A2(n597), .B1(\entry[3][7] ), .B2(n598), 
        .ZN(n652) );
  AOI22D0 U661 ( .A1(\entry[0][7] ), .A2(n599), .B1(\entry[5][7] ), .B2(n600), 
        .ZN(n651) );
  AOI22D0 U662 ( .A1(\entry[1][7] ), .A2(n601), .B1(\entry[7][7] ), .B2(n602), 
        .ZN(n650) );
  AOI22D0 U663 ( .A1(\entry[6][7] ), .A2(n603), .B1(\entry[4][7] ), .B2(n604), 
        .ZN(n649) );
  ND4D0 U664 ( .A1(n653), .A2(n654), .A3(n655), .A4(n656), .ZN(N112) );
  AOI22D0 U665 ( .A1(\entry[2][6] ), .A2(n597), .B1(\entry[3][6] ), .B2(n598), 
        .ZN(n656) );
  AOI22D0 U666 ( .A1(\entry[0][6] ), .A2(n599), .B1(\entry[5][6] ), .B2(n600), 
        .ZN(n655) );
  AOI22D0 U667 ( .A1(\entry[1][6] ), .A2(n601), .B1(\entry[7][6] ), .B2(n602), 
        .ZN(n654) );
  AOI22D0 U668 ( .A1(\entry[6][6] ), .A2(n603), .B1(\entry[4][6] ), .B2(n604), 
        .ZN(n653) );
  ND4D0 U669 ( .A1(n657), .A2(n658), .A3(n659), .A4(n660), .ZN(N111) );
  AOI22D0 U670 ( .A1(\entry[2][5] ), .A2(n597), .B1(\entry[3][5] ), .B2(n598), 
        .ZN(n660) );
  AOI22D0 U671 ( .A1(\entry[0][5] ), .A2(n599), .B1(\entry[5][5] ), .B2(n600), 
        .ZN(n659) );
  AOI22D0 U672 ( .A1(\entry[1][5] ), .A2(n601), .B1(\entry[7][5] ), .B2(n602), 
        .ZN(n658) );
  AOI22D0 U673 ( .A1(\entry[6][5] ), .A2(n603), .B1(\entry[4][5] ), .B2(n604), 
        .ZN(n657) );
  ND4D0 U674 ( .A1(n661), .A2(n662), .A3(n663), .A4(n664), .ZN(N110) );
  AOI22D0 U675 ( .A1(\entry[2][4] ), .A2(n597), .B1(\entry[3][4] ), .B2(n598), 
        .ZN(n664) );
  AOI22D0 U676 ( .A1(\entry[0][4] ), .A2(n599), .B1(\entry[5][4] ), .B2(n600), 
        .ZN(n663) );
  AOI22D0 U677 ( .A1(\entry[1][4] ), .A2(n601), .B1(\entry[7][4] ), .B2(n602), 
        .ZN(n662) );
  AOI22D0 U678 ( .A1(\entry[6][4] ), .A2(n603), .B1(\entry[4][4] ), .B2(n604), 
        .ZN(n661) );
  ND4D0 U679 ( .A1(n665), .A2(n666), .A3(n667), .A4(n668), .ZN(N109) );
  AOI22D0 U680 ( .A1(\entry[2][3] ), .A2(n597), .B1(\entry[3][3] ), .B2(n598), 
        .ZN(n668) );
  AOI22D0 U681 ( .A1(\entry[0][3] ), .A2(n599), .B1(\entry[5][3] ), .B2(n600), 
        .ZN(n667) );
  AOI22D0 U682 ( .A1(\entry[1][3] ), .A2(n601), .B1(\entry[7][3] ), .B2(n602), 
        .ZN(n666) );
  AOI22D0 U683 ( .A1(\entry[6][3] ), .A2(n603), .B1(\entry[4][3] ), .B2(n604), 
        .ZN(n665) );
  ND4D0 U684 ( .A1(n669), .A2(n670), .A3(n671), .A4(n672), .ZN(N108) );
  AOI22D0 U685 ( .A1(\entry[2][2] ), .A2(n597), .B1(\entry[3][2] ), .B2(n598), 
        .ZN(n672) );
  AOI22D0 U686 ( .A1(\entry[0][2] ), .A2(n599), .B1(\entry[5][2] ), .B2(n600), 
        .ZN(n671) );
  AOI22D0 U687 ( .A1(\entry[1][2] ), .A2(n601), .B1(\entry[7][2] ), .B2(n602), 
        .ZN(n670) );
  AOI22D0 U688 ( .A1(\entry[6][2] ), .A2(n603), .B1(\entry[4][2] ), .B2(n604), 
        .ZN(n669) );
  ND4D0 U689 ( .A1(n673), .A2(n674), .A3(n675), .A4(n676), .ZN(N107) );
  AOI22D0 U690 ( .A1(\entry[2][1] ), .A2(n597), .B1(\entry[3][1] ), .B2(n598), 
        .ZN(n676) );
  AOI22D0 U691 ( .A1(\entry[0][1] ), .A2(n599), .B1(\entry[5][1] ), .B2(n600), 
        .ZN(n675) );
  AOI22D0 U692 ( .A1(\entry[1][1] ), .A2(n601), .B1(\entry[7][1] ), .B2(n602), 
        .ZN(n674) );
  AOI22D0 U693 ( .A1(\entry[6][1] ), .A2(n603), .B1(\entry[4][1] ), .B2(n604), 
        .ZN(n673) );
  ND4D0 U694 ( .A1(n677), .A2(n678), .A3(n679), .A4(n680), .ZN(N106) );
  AOI22D0 U695 ( .A1(\entry[2][0] ), .A2(n597), .B1(\entry[3][0] ), .B2(n598), 
        .ZN(n680) );
  AOI22D0 U696 ( .A1(\entry[0][0] ), .A2(n599), .B1(\entry[5][0] ), .B2(n600), 
        .ZN(n679) );
  AOI22D0 U697 ( .A1(\entry[1][0] ), .A2(n601), .B1(\entry[7][0] ), .B2(n602), 
        .ZN(n678) );
  CKND0 U698 ( .I(n681), .ZN(n602) );
  CKND0 U699 ( .I(n682), .ZN(n601) );
  AOI22D0 U700 ( .A1(\entry[6][0] ), .A2(n603), .B1(\entry[4][0] ), .B2(n604), 
        .ZN(n677) );
  NR4D0 U701 ( .A1(n598), .A2(n597), .A3(n604), .A4(n603), .ZN(n684) );
  CKND0 U702 ( .I(n685), .ZN(n603) );
  IND3D0 U703 ( .A1(n686), .B1(n687), .B2(n688), .ZN(n685) );
  IINR4D0 U704 ( .A1(n689), .A2(n690), .B1(n691), .B2(n692), .ZN(n604) );
  AN2D0 U705 ( .A1(n689), .A2(n692), .Z(n597) );
  CKND0 U706 ( .I(n693), .ZN(n598) );
  IND3D0 U707 ( .A1(n692), .B1(n689), .B2(n691), .ZN(n693) );
  NR2D0 U708 ( .A1(n600), .A2(n599), .ZN(n683) );
  AN2D0 U709 ( .A1(n694), .A2(n695), .Z(n599) );
  AN2D0 U710 ( .A1(n687), .A2(n686), .Z(n600) );
  OAI211D0 U711 ( .A1(n696), .A2(n697), .B(n687), .C(n698), .ZN(n681) );
  NR2D0 U712 ( .A1(n688), .A2(n686), .ZN(n698) );
  CKND2D0 U713 ( .A1(n699), .A2(n700), .ZN(n686) );
  AN4D0 U714 ( .A1(n701), .A2(n702), .A3(n703), .A4(n704), .Z(n700) );
  AOI222D0 U715 ( .A1(\entry[5][22] ), .A2(tag[2]), .B1(\entry[5][20] ), .B2(
        tag[0]), .C1(\entry[5][21] ), .C2(tag[1]), .ZN(n704) );
  AOI222D0 U716 ( .A1(\entry[5][25] ), .A2(tag[5]), .B1(\entry[5][23] ), .B2(
        tag[3]), .C1(\entry[5][24] ), .C2(tag[4]), .ZN(n703) );
  AOI222D0 U717 ( .A1(\entry[5][28] ), .A2(tag[8]), .B1(\entry[5][26] ), .B2(
        tag[6]), .C1(\entry[5][27] ), .C2(tag[7]), .ZN(n702) );
  AOI222D0 U718 ( .A1(\entry[5][31] ), .A2(tag[11]), .B1(\entry[5][29] ), .B2(
        tag[9]), .C1(\entry[5][30] ), .C2(tag[10]), .ZN(n701) );
  AN4D0 U719 ( .A1(n705), .A2(n706), .A3(n707), .A4(n708), .Z(n699) );
  AOI222D0 U720 ( .A1(\entry[5][34] ), .A2(tag[14]), .B1(\entry[5][32] ), .B2(
        tag[12]), .C1(\entry[5][33] ), .C2(tag[13]), .ZN(n708) );
  AOI222D0 U721 ( .A1(\entry[5][37] ), .A2(tag[17]), .B1(\entry[5][35] ), .B2(
        tag[15]), .C1(\entry[5][36] ), .C2(tag[16]), .ZN(n707) );
  AOI222D0 U722 ( .A1(\entry[5][40] ), .A2(tag[20]), .B1(\entry[5][38] ), .B2(
        tag[18]), .C1(\entry[5][39] ), .C2(tag[19]), .ZN(n706) );
  AOI222D0 U723 ( .A1(\entry[5][43] ), .A2(tag[23]), .B1(\entry[5][41] ), .B2(
        tag[21]), .C1(\entry[5][42] ), .C2(tag[22]), .ZN(n705) );
  CKND2D0 U724 ( .A1(n709), .A2(n710), .ZN(n688) );
  AN4D0 U725 ( .A1(n711), .A2(n712), .A3(n713), .A4(n714), .Z(n710) );
  AOI222D0 U726 ( .A1(\entry[6][22] ), .A2(tag[2]), .B1(\entry[6][20] ), .B2(
        tag[0]), .C1(\entry[6][21] ), .C2(tag[1]), .ZN(n714) );
  AOI222D0 U727 ( .A1(\entry[6][25] ), .A2(tag[5]), .B1(\entry[6][23] ), .B2(
        tag[3]), .C1(\entry[6][24] ), .C2(tag[4]), .ZN(n713) );
  AOI222D0 U728 ( .A1(\entry[6][28] ), .A2(tag[8]), .B1(\entry[6][26] ), .B2(
        tag[6]), .C1(\entry[6][27] ), .C2(tag[7]), .ZN(n712) );
  AOI222D0 U729 ( .A1(\entry[6][31] ), .A2(tag[11]), .B1(\entry[6][29] ), .B2(
        tag[9]), .C1(\entry[6][30] ), .C2(tag[10]), .ZN(n711) );
  AN4D0 U730 ( .A1(n715), .A2(n716), .A3(n717), .A4(n718), .Z(n709) );
  AOI222D0 U731 ( .A1(\entry[6][34] ), .A2(tag[14]), .B1(\entry[6][32] ), .B2(
        tag[12]), .C1(\entry[6][33] ), .C2(tag[13]), .ZN(n718) );
  AOI222D0 U732 ( .A1(\entry[6][37] ), .A2(tag[17]), .B1(\entry[6][35] ), .B2(
        tag[15]), .C1(\entry[6][36] ), .C2(tag[16]), .ZN(n717) );
  AOI222D0 U733 ( .A1(\entry[6][40] ), .A2(tag[20]), .B1(\entry[6][38] ), .B2(
        tag[18]), .C1(\entry[6][39] ), .C2(tag[19]), .ZN(n716) );
  AOI222D0 U734 ( .A1(\entry[6][43] ), .A2(tag[23]), .B1(\entry[6][41] ), .B2(
        tag[21]), .C1(\entry[6][42] ), .C2(tag[22]), .ZN(n715) );
  INR4D0 U735 ( .A1(n689), .B1(n691), .B2(n690), .B3(n692), .ZN(n687) );
  CKND2D0 U736 ( .A1(n719), .A2(n720), .ZN(n692) );
  AN4D0 U737 ( .A1(n721), .A2(n722), .A3(n723), .A4(n724), .Z(n720) );
  AOI222D0 U738 ( .A1(\entry[2][22] ), .A2(tag[2]), .B1(\entry[2][20] ), .B2(
        tag[0]), .C1(\entry[2][21] ), .C2(tag[1]), .ZN(n724) );
  AOI222D0 U739 ( .A1(\entry[2][25] ), .A2(tag[5]), .B1(\entry[2][23] ), .B2(
        tag[3]), .C1(\entry[2][24] ), .C2(tag[4]), .ZN(n723) );
  AOI222D0 U740 ( .A1(\entry[2][28] ), .A2(tag[8]), .B1(\entry[2][26] ), .B2(
        tag[6]), .C1(\entry[2][27] ), .C2(tag[7]), .ZN(n722) );
  AOI222D0 U741 ( .A1(\entry[2][31] ), .A2(tag[11]), .B1(\entry[2][29] ), .B2(
        tag[9]), .C1(\entry[2][30] ), .C2(tag[10]), .ZN(n721) );
  AN4D0 U742 ( .A1(n725), .A2(n726), .A3(n727), .A4(n728), .Z(n719) );
  AOI222D0 U743 ( .A1(\entry[2][34] ), .A2(tag[14]), .B1(\entry[2][32] ), .B2(
        tag[12]), .C1(\entry[2][33] ), .C2(tag[13]), .ZN(n728) );
  AOI222D0 U744 ( .A1(\entry[2][37] ), .A2(tag[17]), .B1(\entry[2][35] ), .B2(
        tag[15]), .C1(\entry[2][36] ), .C2(tag[16]), .ZN(n727) );
  AOI222D0 U745 ( .A1(\entry[2][40] ), .A2(tag[20]), .B1(\entry[2][38] ), .B2(
        tag[18]), .C1(\entry[2][39] ), .C2(tag[19]), .ZN(n726) );
  AOI222D0 U746 ( .A1(\entry[2][43] ), .A2(tag[23]), .B1(\entry[2][41] ), .B2(
        tag[21]), .C1(\entry[2][42] ), .C2(tag[22]), .ZN(n725) );
  CKND2D0 U747 ( .A1(n729), .A2(n730), .ZN(n690) );
  AN4D0 U748 ( .A1(n731), .A2(n732), .A3(n733), .A4(n734), .Z(n730) );
  AOI222D0 U749 ( .A1(\entry[4][22] ), .A2(tag[2]), .B1(\entry[4][20] ), .B2(
        tag[0]), .C1(\entry[4][21] ), .C2(tag[1]), .ZN(n734) );
  AOI222D0 U750 ( .A1(\entry[4][25] ), .A2(tag[5]), .B1(\entry[4][23] ), .B2(
        tag[3]), .C1(\entry[4][24] ), .C2(tag[4]), .ZN(n733) );
  AOI222D0 U751 ( .A1(\entry[4][28] ), .A2(tag[8]), .B1(\entry[4][26] ), .B2(
        tag[6]), .C1(\entry[4][27] ), .C2(tag[7]), .ZN(n732) );
  AOI222D0 U752 ( .A1(\entry[4][31] ), .A2(tag[11]), .B1(\entry[4][29] ), .B2(
        tag[9]), .C1(\entry[4][30] ), .C2(tag[10]), .ZN(n731) );
  AN4D0 U753 ( .A1(n735), .A2(n736), .A3(n737), .A4(n738), .Z(n729) );
  AOI222D0 U754 ( .A1(\entry[4][34] ), .A2(tag[14]), .B1(\entry[4][32] ), .B2(
        tag[12]), .C1(\entry[4][33] ), .C2(tag[13]), .ZN(n738) );
  AOI222D0 U755 ( .A1(\entry[4][37] ), .A2(tag[17]), .B1(\entry[4][35] ), .B2(
        tag[15]), .C1(\entry[4][36] ), .C2(tag[16]), .ZN(n737) );
  AOI222D0 U756 ( .A1(\entry[4][40] ), .A2(tag[20]), .B1(\entry[4][38] ), .B2(
        tag[18]), .C1(\entry[4][39] ), .C2(tag[19]), .ZN(n736) );
  AOI222D0 U757 ( .A1(\entry[4][43] ), .A2(tag[23]), .B1(\entry[4][41] ), .B2(
        tag[21]), .C1(\entry[4][42] ), .C2(tag[22]), .ZN(n735) );
  CKND2D0 U758 ( .A1(n739), .A2(n740), .ZN(n691) );
  AN4D0 U759 ( .A1(n741), .A2(n742), .A3(n743), .A4(n744), .Z(n740) );
  AOI222D0 U760 ( .A1(\entry[3][22] ), .A2(tag[2]), .B1(\entry[3][20] ), .B2(
        tag[0]), .C1(\entry[3][21] ), .C2(tag[1]), .ZN(n744) );
  AOI222D0 U761 ( .A1(\entry[3][25] ), .A2(tag[5]), .B1(\entry[3][23] ), .B2(
        tag[3]), .C1(\entry[3][24] ), .C2(tag[4]), .ZN(n743) );
  AOI222D0 U762 ( .A1(\entry[3][28] ), .A2(tag[8]), .B1(\entry[3][26] ), .B2(
        tag[6]), .C1(\entry[3][27] ), .C2(tag[7]), .ZN(n742) );
  AOI222D0 U763 ( .A1(\entry[3][31] ), .A2(tag[11]), .B1(\entry[3][29] ), .B2(
        tag[9]), .C1(\entry[3][30] ), .C2(tag[10]), .ZN(n741) );
  AN4D0 U764 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .Z(n739) );
  AOI222D0 U765 ( .A1(\entry[3][34] ), .A2(tag[14]), .B1(\entry[3][32] ), .B2(
        tag[12]), .C1(\entry[3][33] ), .C2(tag[13]), .ZN(n748) );
  AOI222D0 U766 ( .A1(\entry[3][37] ), .A2(tag[17]), .B1(\entry[3][35] ), .B2(
        tag[15]), .C1(\entry[3][36] ), .C2(tag[16]), .ZN(n747) );
  AOI222D0 U767 ( .A1(\entry[3][40] ), .A2(tag[20]), .B1(\entry[3][38] ), .B2(
        tag[18]), .C1(\entry[3][39] ), .C2(tag[19]), .ZN(n746) );
  AOI222D0 U768 ( .A1(\entry[3][43] ), .A2(tag[23]), .B1(\entry[3][41] ), .B2(
        tag[21]), .C1(\entry[3][42] ), .C2(tag[22]), .ZN(n745) );
  INR3D0 U769 ( .A1(n694), .B1(n695), .B2(n749), .ZN(n689) );
  ND4D0 U770 ( .A1(n750), .A2(n751), .A3(n752), .A4(n753), .ZN(n697) );
  AOI222D0 U771 ( .A1(\entry[7][34] ), .A2(tag[14]), .B1(\entry[7][32] ), .B2(
        tag[12]), .C1(\entry[7][33] ), .C2(tag[13]), .ZN(n753) );
  AOI222D0 U772 ( .A1(\entry[7][37] ), .A2(tag[17]), .B1(\entry[7][35] ), .B2(
        tag[15]), .C1(\entry[7][36] ), .C2(tag[16]), .ZN(n752) );
  AOI222D0 U773 ( .A1(\entry[7][40] ), .A2(tag[20]), .B1(\entry[7][38] ), .B2(
        tag[18]), .C1(\entry[7][39] ), .C2(tag[19]), .ZN(n751) );
  AOI222D0 U774 ( .A1(\entry[7][43] ), .A2(tag[23]), .B1(\entry[7][41] ), .B2(
        tag[21]), .C1(\entry[7][42] ), .C2(tag[22]), .ZN(n750) );
  ND4D0 U775 ( .A1(n754), .A2(n755), .A3(n756), .A4(n757), .ZN(n696) );
  AOI222D0 U776 ( .A1(\entry[7][22] ), .A2(tag[2]), .B1(\entry[7][20] ), .B2(
        tag[0]), .C1(\entry[7][21] ), .C2(tag[1]), .ZN(n757) );
  AOI222D0 U777 ( .A1(\entry[7][25] ), .A2(tag[5]), .B1(\entry[7][23] ), .B2(
        tag[3]), .C1(\entry[7][24] ), .C2(tag[4]), .ZN(n756) );
  AOI222D0 U778 ( .A1(\entry[7][28] ), .A2(tag[8]), .B1(\entry[7][26] ), .B2(
        tag[6]), .C1(\entry[7][27] ), .C2(tag[7]), .ZN(n755) );
  AOI222D0 U779 ( .A1(\entry[7][31] ), .A2(tag[11]), .B1(\entry[7][29] ), .B2(
        tag[9]), .C1(\entry[7][30] ), .C2(tag[10]), .ZN(n754) );
  IND3D0 U780 ( .A1(n695), .B1(n749), .B2(n694), .ZN(n682) );
  NR2D0 U781 ( .A1(rst), .A2(wr), .ZN(n694) );
  CKND2D0 U782 ( .A1(n758), .A2(n759), .ZN(n749) );
  AN4D0 U783 ( .A1(n760), .A2(n761), .A3(n762), .A4(n763), .Z(n759) );
  AOI222D0 U784 ( .A1(\entry[1][22] ), .A2(tag[2]), .B1(\entry[1][20] ), .B2(
        tag[0]), .C1(\entry[1][21] ), .C2(tag[1]), .ZN(n763) );
  AOI222D0 U785 ( .A1(\entry[1][25] ), .A2(tag[5]), .B1(\entry[1][23] ), .B2(
        tag[3]), .C1(\entry[1][24] ), .C2(tag[4]), .ZN(n762) );
  AOI222D0 U786 ( .A1(\entry[1][28] ), .A2(tag[8]), .B1(\entry[1][26] ), .B2(
        tag[6]), .C1(\entry[1][27] ), .C2(tag[7]), .ZN(n761) );
  AOI222D0 U787 ( .A1(\entry[1][31] ), .A2(tag[11]), .B1(\entry[1][29] ), .B2(
        tag[9]), .C1(\entry[1][30] ), .C2(tag[10]), .ZN(n760) );
  AN4D0 U788 ( .A1(n764), .A2(n765), .A3(n766), .A4(n767), .Z(n758) );
  AOI222D0 U789 ( .A1(\entry[1][34] ), .A2(tag[14]), .B1(\entry[1][32] ), .B2(
        tag[12]), .C1(\entry[1][33] ), .C2(tag[13]), .ZN(n767) );
  AOI222D0 U790 ( .A1(\entry[1][37] ), .A2(tag[17]), .B1(\entry[1][35] ), .B2(
        tag[15]), .C1(\entry[1][36] ), .C2(tag[16]), .ZN(n766) );
  AOI222D0 U791 ( .A1(\entry[1][40] ), .A2(tag[20]), .B1(\entry[1][38] ), .B2(
        tag[18]), .C1(\entry[1][39] ), .C2(tag[19]), .ZN(n765) );
  AOI222D0 U792 ( .A1(\entry[1][43] ), .A2(tag[23]), .B1(\entry[1][41] ), .B2(
        tag[21]), .C1(\entry[1][42] ), .C2(tag[22]), .ZN(n764) );
  CKND2D0 U793 ( .A1(n768), .A2(n769), .ZN(n695) );
  AN4D0 U794 ( .A1(n770), .A2(n771), .A3(n772), .A4(n773), .Z(n769) );
  AOI222D0 U795 ( .A1(\entry[0][22] ), .A2(tag[2]), .B1(\entry[0][20] ), .B2(
        tag[0]), .C1(\entry[0][21] ), .C2(tag[1]), .ZN(n773) );
  AOI222D0 U796 ( .A1(\entry[0][25] ), .A2(tag[5]), .B1(\entry[0][23] ), .B2(
        tag[3]), .C1(\entry[0][24] ), .C2(tag[4]), .ZN(n772) );
  AOI222D0 U797 ( .A1(\entry[0][28] ), .A2(tag[8]), .B1(\entry[0][26] ), .B2(
        tag[6]), .C1(\entry[0][27] ), .C2(tag[7]), .ZN(n771) );
  AOI222D0 U798 ( .A1(\entry[0][31] ), .A2(tag[11]), .B1(\entry[0][29] ), .B2(
        tag[9]), .C1(\entry[0][30] ), .C2(tag[10]), .ZN(n770) );
  AN4D0 U799 ( .A1(n774), .A2(n775), .A3(n776), .A4(n777), .Z(n768) );
  AOI222D0 U800 ( .A1(\entry[0][34] ), .A2(tag[14]), .B1(\entry[0][32] ), .B2(
        tag[12]), .C1(\entry[0][33] ), .C2(tag[13]), .ZN(n777) );
  AOI222D0 U801 ( .A1(\entry[0][37] ), .A2(tag[17]), .B1(\entry[0][35] ), .B2(
        tag[15]), .C1(\entry[0][36] ), .C2(tag[16]), .ZN(n776) );
  AOI222D0 U802 ( .A1(\entry[0][40] ), .A2(tag[20]), .B1(\entry[0][38] ), .B2(
        tag[18]), .C1(\entry[0][39] ), .C2(tag[19]), .ZN(n775) );
  AOI222D0 U803 ( .A1(\entry[0][43] ), .A2(tag[23]), .B1(\entry[0][41] ), .B2(
        tag[21]), .C1(\entry[0][42] ), .C2(tag[22]), .ZN(n774) );
  OAI211D0 U804 ( .A1(n588), .A2(n778), .B(n585), .C(n590), .ZN(N104) );
  CKND2D0 U805 ( .A1(count[2]), .A2(N102), .ZN(n585) );
  CKND2D0 U806 ( .A1(n780), .A2(n586), .ZN(n778) );
  OAI21D0 U807 ( .A1(n591), .A2(n586), .B(n589), .ZN(N103) );
  ND3D0 U808 ( .A1(n780), .A2(n586), .A3(count[0]), .ZN(n589) );
  CKND0 U809 ( .I(count[1]), .ZN(n586) );
  CKND0 U810 ( .I(N102), .ZN(n591) );
  NR2D0 U811 ( .A1(n592), .A2(count[0]), .ZN(N102) );
  CKND2D0 U812 ( .A1(n587), .A2(n592), .ZN(N101) );
  ND3D0 U813 ( .A1(count[1]), .A2(n780), .A3(count[0]), .ZN(n779) );
  CKND0 U814 ( .I(n592), .ZN(n780) );
  CKND2D0 U815 ( .A1(wr), .A2(n587), .ZN(n592) );
  CKND0 U816 ( .I(rst), .ZN(n587) );
  CKND0 U817 ( .I(count[2]), .ZN(n588) );
endmodule

