
module activationFunction ( clk, rst, wr, index, val, store_val, boundary_val, 
        en, out_coef, out_bias );
  input [3:0] index;
  input [15:0] val;
  input [31:0] store_val;
  input [15:0] boundary_val;
  output [15:0] out_coef;
  output [15:0] out_bias;
  input clk, rst, wr, en;
  wire   \entry[15][31] , \entry[15][30] , \entry[15][29] , \entry[15][28] ,
         \entry[15][27] , \entry[15][26] , \entry[15][25] , \entry[15][24] ,
         \entry[15][23] , \entry[15][22] , \entry[15][21] , \entry[15][20] ,
         \entry[15][19] , \entry[15][18] , \entry[15][17] , \entry[15][16] ,
         \entry[15][15] , \entry[15][14] , \entry[15][13] , \entry[15][12] ,
         \entry[15][11] , \entry[15][10] , \entry[15][9] , \entry[15][8] ,
         \entry[15][7] , \entry[15][6] , \entry[15][5] , \entry[15][4] ,
         \entry[15][3] , \entry[15][2] , \entry[15][1] , \entry[15][0] ,
         \entry[14][31] , \entry[14][30] , \entry[14][29] , \entry[14][28] ,
         \entry[14][27] , \entry[14][26] , \entry[14][25] , \entry[14][24] ,
         \entry[14][23] , \entry[14][22] , \entry[14][21] , \entry[14][20] ,
         \entry[14][19] , \entry[14][18] , \entry[14][17] , \entry[14][16] ,
         \entry[14][15] , \entry[14][14] , \entry[14][13] , \entry[14][12] ,
         \entry[14][11] , \entry[14][10] , \entry[14][9] , \entry[14][8] ,
         \entry[14][7] , \entry[14][6] , \entry[14][5] , \entry[14][4] ,
         \entry[14][3] , \entry[14][2] , \entry[14][1] , \entry[14][0] ,
         \entry[13][31] , \entry[13][30] , \entry[13][29] , \entry[13][28] ,
         \entry[13][27] , \entry[13][26] , \entry[13][25] , \entry[13][24] ,
         \entry[13][23] , \entry[13][22] , \entry[13][21] , \entry[13][20] ,
         \entry[13][19] , \entry[13][18] , \entry[13][17] , \entry[13][16] ,
         \entry[13][15] , \entry[13][14] , \entry[13][13] , \entry[13][12] ,
         \entry[13][11] , \entry[13][10] , \entry[13][9] , \entry[13][8] ,
         \entry[13][7] , \entry[13][6] , \entry[13][5] , \entry[13][4] ,
         \entry[13][3] , \entry[13][2] , \entry[13][1] , \entry[13][0] ,
         \entry[12][31] , \entry[12][30] , \entry[12][29] , \entry[12][28] ,
         \entry[12][27] , \entry[12][26] , \entry[12][25] , \entry[12][24] ,
         \entry[12][23] , \entry[12][22] , \entry[12][21] , \entry[12][20] ,
         \entry[12][19] , \entry[12][18] , \entry[12][17] , \entry[12][16] ,
         \entry[12][15] , \entry[12][14] , \entry[12][13] , \entry[12][12] ,
         \entry[12][11] , \entry[12][10] , \entry[12][9] , \entry[12][8] ,
         \entry[12][7] , \entry[12][6] , \entry[12][5] , \entry[12][4] ,
         \entry[12][3] , \entry[12][2] , \entry[12][1] , \entry[12][0] ,
         \entry[11][31] , \entry[11][30] , \entry[11][29] , \entry[11][28] ,
         \entry[11][27] , \entry[11][26] , \entry[11][25] , \entry[11][24] ,
         \entry[11][23] , \entry[11][22] , \entry[11][21] , \entry[11][20] ,
         \entry[11][19] , \entry[11][18] , \entry[11][17] , \entry[11][16] ,
         \entry[11][15] , \entry[11][14] , \entry[11][13] , \entry[11][12] ,
         \entry[11][11] , \entry[11][10] , \entry[11][9] , \entry[11][8] ,
         \entry[11][7] , \entry[11][6] , \entry[11][5] , \entry[11][4] ,
         \entry[11][3] , \entry[11][2] , \entry[11][1] , \entry[11][0] ,
         \entry[10][31] , \entry[10][30] , \entry[10][29] , \entry[10][28] ,
         \entry[10][27] , \entry[10][26] , \entry[10][25] , \entry[10][24] ,
         \entry[10][23] , \entry[10][22] , \entry[10][21] , \entry[10][20] ,
         \entry[10][19] , \entry[10][18] , \entry[10][17] , \entry[10][16] ,
         \entry[10][15] , \entry[10][14] , \entry[10][13] , \entry[10][12] ,
         \entry[10][11] , \entry[10][10] , \entry[10][9] , \entry[10][8] ,
         \entry[10][7] , \entry[10][6] , \entry[10][5] , \entry[10][4] ,
         \entry[10][3] , \entry[10][2] , \entry[10][1] , \entry[10][0] ,
         \entry[9][31] , \entry[9][30] , \entry[9][29] , \entry[9][28] ,
         \entry[9][27] , \entry[9][26] , \entry[9][25] , \entry[9][24] ,
         \entry[9][23] , \entry[9][22] , \entry[9][21] , \entry[9][20] ,
         \entry[9][19] , \entry[9][18] , \entry[9][17] , \entry[9][16] ,
         \entry[9][15] , \entry[9][14] , \entry[9][13] , \entry[9][12] ,
         \entry[9][11] , \entry[9][10] , \entry[9][9] , \entry[9][8] ,
         \entry[9][7] , \entry[9][6] , \entry[9][5] , \entry[9][4] ,
         \entry[9][3] , \entry[9][2] , \entry[9][1] , \entry[9][0] ,
         \entry[8][31] , \entry[8][30] , \entry[8][29] , \entry[8][28] ,
         \entry[8][27] , \entry[8][26] , \entry[8][25] , \entry[8][24] ,
         \entry[8][23] , \entry[8][22] , \entry[8][21] , \entry[8][20] ,
         \entry[8][19] , \entry[8][18] , \entry[8][17] , \entry[8][16] ,
         \entry[8][15] , \entry[8][14] , \entry[8][13] , \entry[8][12] ,
         \entry[8][11] , \entry[8][10] , \entry[8][9] , \entry[8][8] ,
         \entry[8][7] , \entry[8][6] , \entry[8][5] , \entry[8][4] ,
         \entry[8][3] , \entry[8][2] , \entry[8][1] , \entry[8][0] ,
         \entry[7][31] , \entry[7][30] , \entry[7][29] , \entry[7][28] ,
         \entry[7][27] , \entry[7][26] , \entry[7][25] , \entry[7][24] ,
         \entry[7][23] , \entry[7][22] , \entry[7][21] , \entry[7][20] ,
         \entry[7][19] , \entry[7][18] , \entry[7][17] , \entry[7][16] ,
         \entry[7][15] , \entry[7][14] , \entry[7][13] , \entry[7][12] ,
         \entry[7][11] , \entry[7][10] , \entry[7][9] , \entry[7][8] ,
         \entry[7][7] , \entry[7][6] , \entry[7][5] , \entry[7][4] ,
         \entry[7][3] , \entry[7][2] , \entry[7][1] , \entry[7][0] ,
         \entry[6][31] , \entry[6][30] , \entry[6][29] , \entry[6][28] ,
         \entry[6][27] , \entry[6][26] , \entry[6][25] , \entry[6][24] ,
         \entry[6][23] , \entry[6][22] , \entry[6][21] , \entry[6][20] ,
         \entry[6][19] , \entry[6][18] , \entry[6][17] , \entry[6][16] ,
         \entry[6][15] , \entry[6][14] , \entry[6][13] , \entry[6][12] ,
         \entry[6][11] , \entry[6][10] , \entry[6][9] , \entry[6][8] ,
         \entry[6][7] , \entry[6][6] , \entry[6][5] , \entry[6][4] ,
         \entry[6][3] , \entry[6][2] , \entry[6][1] , \entry[6][0] ,
         \entry[5][31] , \entry[5][30] , \entry[5][29] , \entry[5][28] ,
         \entry[5][27] , \entry[5][26] , \entry[5][25] , \entry[5][24] ,
         \entry[5][23] , \entry[5][22] , \entry[5][21] , \entry[5][20] ,
         \entry[5][19] , \entry[5][18] , \entry[5][17] , \entry[5][16] ,
         \entry[5][15] , \entry[5][14] , \entry[5][13] , \entry[5][12] ,
         \entry[5][11] , \entry[5][10] , \entry[5][9] , \entry[5][8] ,
         \entry[5][7] , \entry[5][6] , \entry[5][5] , \entry[5][4] ,
         \entry[5][3] , \entry[5][2] , \entry[5][1] , \entry[5][0] ,
         \entry[4][31] , \entry[4][30] , \entry[4][29] , \entry[4][28] ,
         \entry[4][27] , \entry[4][26] , \entry[4][25] , \entry[4][24] ,
         \entry[4][23] , \entry[4][22] , \entry[4][21] , \entry[4][20] ,
         \entry[4][19] , \entry[4][18] , \entry[4][17] , \entry[4][16] ,
         \entry[4][15] , \entry[4][14] , \entry[4][13] , \entry[4][12] ,
         \entry[4][11] , \entry[4][10] , \entry[4][9] , \entry[4][8] ,
         \entry[4][7] , \entry[4][6] , \entry[4][5] , \entry[4][4] ,
         \entry[4][3] , \entry[4][2] , \entry[4][1] , \entry[4][0] ,
         \entry[3][31] , \entry[3][30] , \entry[3][29] , \entry[3][28] ,
         \entry[3][27] , \entry[3][26] , \entry[3][25] , \entry[3][24] ,
         \entry[3][23] , \entry[3][22] , \entry[3][21] , \entry[3][20] ,
         \entry[3][19] , \entry[3][18] , \entry[3][17] , \entry[3][16] ,
         \entry[3][15] , \entry[3][14] , \entry[3][13] , \entry[3][12] ,
         \entry[3][11] , \entry[3][10] , \entry[3][9] , \entry[3][8] ,
         \entry[3][7] , \entry[3][6] , \entry[3][5] , \entry[3][4] ,
         \entry[3][3] , \entry[3][2] , \entry[3][1] , \entry[3][0] ,
         \entry[2][31] , \entry[2][30] , \entry[2][29] , \entry[2][28] ,
         \entry[2][27] , \entry[2][26] , \entry[2][25] , \entry[2][24] ,
         \entry[2][23] , \entry[2][22] , \entry[2][21] , \entry[2][20] ,
         \entry[2][19] , \entry[2][18] , \entry[2][17] , \entry[2][16] ,
         \entry[2][15] , \entry[2][14] , \entry[2][13] , \entry[2][12] ,
         \entry[2][11] , \entry[2][10] , \entry[2][9] , \entry[2][8] ,
         \entry[2][7] , \entry[2][6] , \entry[2][5] , \entry[2][4] ,
         \entry[2][3] , \entry[2][2] , \entry[2][1] , \entry[2][0] ,
         \entry[1][31] , \entry[1][30] , \entry[1][29] , \entry[1][28] ,
         \entry[1][27] , \entry[1][26] , \entry[1][25] , \entry[1][24] ,
         \entry[1][23] , \entry[1][22] , \entry[1][21] , \entry[1][20] ,
         \entry[1][19] , \entry[1][18] , \entry[1][17] , \entry[1][16] ,
         \entry[1][15] , \entry[1][14] , \entry[1][13] , \entry[1][12] ,
         \entry[1][11] , \entry[1][10] , \entry[1][9] , \entry[1][8] ,
         \entry[1][7] , \entry[1][6] , \entry[1][5] , \entry[1][4] ,
         \entry[1][3] , \entry[1][2] , \entry[1][1] , \entry[1][0] ,
         \entry[0][31] , \entry[0][30] , \entry[0][29] , \entry[0][28] ,
         \entry[0][27] , \entry[0][26] , \entry[0][25] , \entry[0][24] ,
         \entry[0][23] , \entry[0][22] , \entry[0][21] , \entry[0][20] ,
         \entry[0][19] , \entry[0][18] , \entry[0][17] , \entry[0][16] ,
         \entry[0][15] , \entry[0][14] , \entry[0][13] , \entry[0][12] ,
         \entry[0][11] , \entry[0][10] , \entry[0][9] , \entry[0][8] ,
         \entry[0][7] , \entry[0][6] , \entry[0][5] , \entry[0][4] ,
         \entry[0][3] , \entry[0][2] , \entry[0][1] , \entry[0][0] , N10284,
         N10285, N10286, N10287, N10288, N10289, N10290, N10291, N10292,
         N10293, N10294, N10295, N10296, N10297, N10298, N10299, N10301,
         N10302, N10303, N10304, N10305, N10306, N10307, N10308, N10309,
         N10310, N10311, N10312, N10313, N10314, N10315, N10316, N10317,
         N10318, N10319, N10320, N10321, N10322, N10323, N10324, N10325,
         N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333,
         N10334, N10335, N10336, N10337, N10338, N10339, N10340, N10341,
         N10342, N10343, N10344, N10345, N10346, N10347, N10348, N10349,
         N10350, N10351, N10352, N10353, N10354, N10355, N10356, N10357,
         N10358, N10359, N10360, N10361, N10362, N10363, N10364, N10366, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2463, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343;

  LHD1 \boundary_flags_reg[14][0]  ( .E(n2463), .D(n2463), .QN(n2182) );
  LHD1 \boundary_flags_reg[14][1]  ( .E(n2463), .D(n2463), .QN(n2181) );
  LHD1 \boundary_flags_reg[12][0]  ( .E(n2463), .D(n2463), .QN(n2186) );
  LHD1 \boundary_flags_reg[12][1]  ( .E(n2463), .D(n2463), .QN(n2185) );
  LHD1 \boundary_flags_reg[10][0]  ( .E(n2463), .D(n2463), .QN(n2194) );
  LHD1 \boundary_flags_reg[10][1]  ( .E(n2463), .D(n2463), .QN(n2193) );
  LHD1 \boundary_flags_reg[8][0]  ( .E(n2463), .D(n2463), .QN(n2190) );
  LHD1 \boundary_flags_reg[8][1]  ( .E(n2463), .D(n2463), .QN(n2189) );
  LHD1 \boundary_flags_reg[6][0]  ( .E(n2463), .D(n2463), .QN(n2198) );
  LHD1 \boundary_flags_reg[6][1]  ( .E(n2463), .D(n2463), .QN(n2197) );
  LHD1 \boundary_flags_reg[4][0]  ( .E(n2463), .D(n2463), .QN(n2202) );
  LHD1 \boundary_flags_reg[4][1]  ( .E(n2463), .D(n2463), .QN(n2201) );
  LHD1 \boundary_flags_reg[2][0]  ( .E(n2463), .D(n2463), .QN(n2206) );
  LHD1 \boundary_flags_reg[2][1]  ( .E(n2463), .D(n2463), .QN(n2205) );
  LHD1 \boundary_flags_reg[0][0]  ( .E(n2463), .D(n2463), .QN(n3343) );
  LHD1 \boundary_flags_reg[0][1]  ( .E(n2463), .D(n2463), .QN(n3342) );
  LHD1 \boundary_flags_reg[15][0]  ( .E(n2463), .D(n2463), .QN(n3340) );
  LHD1 \boundary_flags_reg[15][1]  ( .E(n2463), .D(n2463), .QN(n3341) );
  LHD1 \boundary_flags_reg[13][0]  ( .E(n2463), .D(n2463), .QN(n2184) );
  LHD1 \boundary_flags_reg[13][1]  ( .E(n2463), .D(n2463), .QN(n2183) );
  LHD1 \boundary_flags_reg[11][0]  ( .E(n2463), .D(n2463), .QN(n2188) );
  LHD1 \boundary_flags_reg[11][1]  ( .E(n2463), .D(n2463), .QN(n2187) );
  LHD1 \boundary_flags_reg[9][0]  ( .E(n2463), .D(n2463), .QN(n2192) );
  LHD1 \boundary_flags_reg[9][1]  ( .E(n2463), .D(n2463), .QN(n2191) );
  LHD1 \boundary_flags_reg[7][0]  ( .E(n2463), .D(n2463), .QN(n2196) );
  LHD1 \boundary_flags_reg[7][1]  ( .E(n2463), .D(n2463), .QN(n2195) );
  LHD1 \boundary_flags_reg[5][0]  ( .E(n2463), .D(n2463), .QN(n2200) );
  LHD1 \boundary_flags_reg[5][1]  ( .E(n2463), .D(n2463), .QN(n2199) );
  LHD1 \boundary_flags_reg[3][0]  ( .E(n2463), .D(n2463), .QN(n2208) );
  LHD1 \boundary_flags_reg[3][1]  ( .E(n2463), .D(n2463), .QN(n2207) );
  LHD1 \boundary_flags_reg[1][0]  ( .E(n2463), .D(n2463), .QN(n2204) );
  LHD1 \boundary_flags_reg[1][1]  ( .E(n2463), .D(n2463), .QN(n2203) );
  EDFQD2 \out_coef_reg[15]  ( .D(N10299), .E(N10366), .CP(clk), .Q(
        out_coef[15]) );
  EDFQD2 \out_coef_reg[14]  ( .D(N10298), .E(N10366), .CP(clk), .Q(
        out_coef[14]) );
  EDFQD2 \out_coef_reg[13]  ( .D(N10297), .E(N10366), .CP(clk), .Q(
        out_coef[13]) );
  EDFQD2 \out_coef_reg[12]  ( .D(N10296), .E(N10366), .CP(clk), .Q(
        out_coef[12]) );
  EDFQD2 \out_coef_reg[11]  ( .D(N10295), .E(N10366), .CP(clk), .Q(
        out_coef[11]) );
  EDFQD2 \out_coef_reg[10]  ( .D(N10294), .E(N10366), .CP(clk), .Q(
        out_coef[10]) );
  EDFQD2 \out_coef_reg[9]  ( .D(N10293), .E(N10366), .CP(clk), .Q(out_coef[9])
         );
  EDFQD2 \out_coef_reg[8]  ( .D(N10292), .E(N10366), .CP(clk), .Q(out_coef[8])
         );
  EDFQD2 \out_coef_reg[7]  ( .D(N10291), .E(N10366), .CP(clk), .Q(out_coef[7])
         );
  EDFQD2 \out_coef_reg[6]  ( .D(N10290), .E(N10366), .CP(clk), .Q(out_coef[6])
         );
  EDFQD2 \out_coef_reg[5]  ( .D(N10289), .E(N10366), .CP(clk), .Q(out_coef[5])
         );
  EDFQD2 \out_coef_reg[4]  ( .D(N10288), .E(N10366), .CP(clk), .Q(out_coef[4])
         );
  EDFQD2 \out_coef_reg[3]  ( .D(N10287), .E(N10366), .CP(clk), .Q(out_coef[3])
         );
  EDFQD2 \out_coef_reg[2]  ( .D(N10286), .E(N10366), .CP(clk), .Q(out_coef[2])
         );
  EDFQD2 \out_coef_reg[1]  ( .D(N10285), .E(N10366), .CP(clk), .Q(out_coef[1])
         );
  EDFQD2 \out_coef_reg[0]  ( .D(N10284), .E(N10366), .CP(clk), .Q(out_coef[0])
         );
  EDFQD2 \out_bias_reg[15]  ( .D(N10316), .E(N10366), .CP(clk), .Q(
        out_bias[15]) );
  EDFQD2 \out_bias_reg[14]  ( .D(N10315), .E(N10366), .CP(clk), .Q(
        out_bias[14]) );
  EDFQD2 \out_bias_reg[13]  ( .D(N10314), .E(N10366), .CP(clk), .Q(
        out_bias[13]) );
  EDFQD2 \out_bias_reg[12]  ( .D(N10313), .E(N10366), .CP(clk), .Q(
        out_bias[12]) );
  EDFQD2 \out_bias_reg[11]  ( .D(N10312), .E(N10366), .CP(clk), .Q(
        out_bias[11]) );
  EDFQD2 \out_bias_reg[10]  ( .D(N10311), .E(N10366), .CP(clk), .Q(
        out_bias[10]) );
  EDFQD2 \out_bias_reg[9]  ( .D(N10310), .E(N10366), .CP(clk), .Q(out_bias[9])
         );
  EDFQD2 \out_bias_reg[8]  ( .D(N10309), .E(N10366), .CP(clk), .Q(out_bias[8])
         );
  EDFQD2 \out_bias_reg[7]  ( .D(N10308), .E(N10366), .CP(clk), .Q(out_bias[7])
         );
  EDFQD2 \out_bias_reg[6]  ( .D(N10307), .E(N10366), .CP(clk), .Q(out_bias[6])
         );
  EDFQD2 \out_bias_reg[5]  ( .D(N10306), .E(N10366), .CP(clk), .Q(out_bias[5])
         );
  EDFQD2 \out_bias_reg[4]  ( .D(N10305), .E(N10366), .CP(clk), .Q(out_bias[4])
         );
  EDFQD2 \out_bias_reg[3]  ( .D(N10304), .E(N10366), .CP(clk), .Q(out_bias[3])
         );
  EDFQD2 \out_bias_reg[2]  ( .D(N10303), .E(N10366), .CP(clk), .Q(out_bias[2])
         );
  EDFQD2 \out_bias_reg[1]  ( .D(N10302), .E(N10366), .CP(clk), .Q(out_bias[1])
         );
  EDFQD2 \out_bias_reg[0]  ( .D(N10301), .E(N10366), .CP(clk), .Q(out_bias[0])
         );
  EDFQD1 \entry_reg[15][31]  ( .D(N10348), .E(N10364), .CP(clk), .Q(
        \entry[15][31] ) );
  EDFQD1 \entry_reg[15][30]  ( .D(N10347), .E(N10364), .CP(clk), .Q(
        \entry[15][30] ) );
  EDFQD1 \entry_reg[15][29]  ( .D(N10346), .E(N10364), .CP(clk), .Q(
        \entry[15][29] ) );
  EDFQD1 \entry_reg[15][28]  ( .D(N10345), .E(N10364), .CP(clk), .Q(
        \entry[15][28] ) );
  EDFQD1 \entry_reg[15][27]  ( .D(N10344), .E(N10364), .CP(clk), .Q(
        \entry[15][27] ) );
  EDFQD1 \entry_reg[15][26]  ( .D(N10343), .E(N10364), .CP(clk), .Q(
        \entry[15][26] ) );
  EDFQD1 \entry_reg[15][25]  ( .D(N10342), .E(N10364), .CP(clk), .Q(
        \entry[15][25] ) );
  EDFQD1 \entry_reg[15][24]  ( .D(N10341), .E(N10364), .CP(clk), .Q(
        \entry[15][24] ) );
  EDFQD1 \entry_reg[15][23]  ( .D(N10340), .E(N10364), .CP(clk), .Q(
        \entry[15][23] ) );
  EDFQD1 \entry_reg[15][22]  ( .D(N10339), .E(N10364), .CP(clk), .Q(
        \entry[15][22] ) );
  EDFQD1 \entry_reg[15][21]  ( .D(N10338), .E(N10364), .CP(clk), .Q(
        \entry[15][21] ) );
  EDFQD1 \entry_reg[15][20]  ( .D(N10337), .E(N10364), .CP(clk), .Q(
        \entry[15][20] ) );
  EDFQD1 \entry_reg[15][19]  ( .D(N10336), .E(N10364), .CP(clk), .Q(
        \entry[15][19] ) );
  EDFQD1 \entry_reg[15][18]  ( .D(N10335), .E(N10364), .CP(clk), .Q(
        \entry[15][18] ) );
  EDFQD1 \entry_reg[15][17]  ( .D(N10334), .E(N10364), .CP(clk), .Q(
        \entry[15][17] ) );
  EDFQD1 \entry_reg[15][16]  ( .D(N10333), .E(N10364), .CP(clk), .Q(
        \entry[15][16] ) );
  EDFQD1 \entry_reg[15][15]  ( .D(N10332), .E(N10364), .CP(clk), .Q(
        \entry[15][15] ) );
  EDFQD1 \entry_reg[15][14]  ( .D(N10331), .E(N10364), .CP(clk), .Q(
        \entry[15][14] ) );
  EDFQD1 \entry_reg[15][13]  ( .D(N10330), .E(N10364), .CP(clk), .Q(
        \entry[15][13] ) );
  EDFQD1 \entry_reg[15][12]  ( .D(N10329), .E(N10364), .CP(clk), .Q(
        \entry[15][12] ) );
  EDFQD1 \entry_reg[15][11]  ( .D(N10328), .E(N10364), .CP(clk), .Q(
        \entry[15][11] ) );
  EDFQD1 \entry_reg[15][10]  ( .D(N10327), .E(N10364), .CP(clk), .Q(
        \entry[15][10] ) );
  EDFQD1 \entry_reg[15][9]  ( .D(N10326), .E(N10364), .CP(clk), .Q(
        \entry[15][9] ) );
  EDFQD1 \entry_reg[15][8]  ( .D(N10325), .E(N10364), .CP(clk), .Q(
        \entry[15][8] ) );
  EDFQD1 \entry_reg[15][7]  ( .D(N10324), .E(N10364), .CP(clk), .Q(
        \entry[15][7] ) );
  EDFQD1 \entry_reg[15][6]  ( .D(N10323), .E(N10364), .CP(clk), .Q(
        \entry[15][6] ) );
  EDFQD1 \entry_reg[15][5]  ( .D(N10322), .E(N10364), .CP(clk), .Q(
        \entry[15][5] ) );
  EDFQD1 \entry_reg[15][4]  ( .D(N10321), .E(N10364), .CP(clk), .Q(
        \entry[15][4] ) );
  EDFQD1 \entry_reg[15][3]  ( .D(N10320), .E(N10364), .CP(clk), .Q(
        \entry[15][3] ) );
  EDFQD1 \entry_reg[15][2]  ( .D(N10319), .E(N10364), .CP(clk), .Q(
        \entry[15][2] ) );
  EDFQD1 \entry_reg[15][1]  ( .D(N10318), .E(N10364), .CP(clk), .Q(
        \entry[15][1] ) );
  EDFQD1 \entry_reg[15][0]  ( .D(N10317), .E(N10364), .CP(clk), .Q(
        \entry[15][0] ) );
  EDFQD1 \entry_reg[14][31]  ( .D(N10348), .E(N10363), .CP(clk), .Q(
        \entry[14][31] ) );
  EDFQD1 \entry_reg[14][30]  ( .D(N10347), .E(N10363), .CP(clk), .Q(
        \entry[14][30] ) );
  EDFQD1 \entry_reg[14][29]  ( .D(N10346), .E(N10363), .CP(clk), .Q(
        \entry[14][29] ) );
  EDFQD1 \entry_reg[14][28]  ( .D(N10345), .E(N10363), .CP(clk), .Q(
        \entry[14][28] ) );
  EDFQD1 \entry_reg[14][27]  ( .D(N10344), .E(N10363), .CP(clk), .Q(
        \entry[14][27] ) );
  EDFQD1 \entry_reg[14][26]  ( .D(N10343), .E(N10363), .CP(clk), .Q(
        \entry[14][26] ) );
  EDFQD1 \entry_reg[14][25]  ( .D(N10342), .E(N10363), .CP(clk), .Q(
        \entry[14][25] ) );
  EDFQD1 \entry_reg[14][24]  ( .D(N10341), .E(N10363), .CP(clk), .Q(
        \entry[14][24] ) );
  EDFQD1 \entry_reg[14][23]  ( .D(N10340), .E(N10363), .CP(clk), .Q(
        \entry[14][23] ) );
  EDFQD1 \entry_reg[14][22]  ( .D(N10339), .E(N10363), .CP(clk), .Q(
        \entry[14][22] ) );
  EDFQD1 \entry_reg[14][21]  ( .D(N10338), .E(N10363), .CP(clk), .Q(
        \entry[14][21] ) );
  EDFQD1 \entry_reg[14][20]  ( .D(N10337), .E(N10363), .CP(clk), .Q(
        \entry[14][20] ) );
  EDFQD1 \entry_reg[14][19]  ( .D(N10336), .E(N10363), .CP(clk), .Q(
        \entry[14][19] ) );
  EDFQD1 \entry_reg[14][18]  ( .D(N10335), .E(N10363), .CP(clk), .Q(
        \entry[14][18] ) );
  EDFQD1 \entry_reg[14][17]  ( .D(N10334), .E(N10363), .CP(clk), .Q(
        \entry[14][17] ) );
  EDFQD1 \entry_reg[14][16]  ( .D(N10333), .E(N10363), .CP(clk), .Q(
        \entry[14][16] ) );
  EDFQD1 \entry_reg[14][15]  ( .D(N10332), .E(N10363), .CP(clk), .Q(
        \entry[14][15] ) );
  EDFQD1 \entry_reg[14][14]  ( .D(N10331), .E(N10363), .CP(clk), .Q(
        \entry[14][14] ) );
  EDFQD1 \entry_reg[14][13]  ( .D(N10330), .E(N10363), .CP(clk), .Q(
        \entry[14][13] ) );
  EDFQD1 \entry_reg[14][12]  ( .D(N10329), .E(N10363), .CP(clk), .Q(
        \entry[14][12] ) );
  EDFQD1 \entry_reg[14][11]  ( .D(N10328), .E(N10363), .CP(clk), .Q(
        \entry[14][11] ) );
  EDFQD1 \entry_reg[14][10]  ( .D(N10327), .E(N10363), .CP(clk), .Q(
        \entry[14][10] ) );
  EDFQD1 \entry_reg[14][9]  ( .D(N10326), .E(N10363), .CP(clk), .Q(
        \entry[14][9] ) );
  EDFQD1 \entry_reg[14][8]  ( .D(N10325), .E(N10363), .CP(clk), .Q(
        \entry[14][8] ) );
  EDFQD1 \entry_reg[14][7]  ( .D(N10324), .E(N10363), .CP(clk), .Q(
        \entry[14][7] ) );
  EDFQD1 \entry_reg[14][6]  ( .D(N10323), .E(N10363), .CP(clk), .Q(
        \entry[14][6] ) );
  EDFQD1 \entry_reg[14][5]  ( .D(N10322), .E(N10363), .CP(clk), .Q(
        \entry[14][5] ) );
  EDFQD1 \entry_reg[14][4]  ( .D(N10321), .E(N10363), .CP(clk), .Q(
        \entry[14][4] ) );
  EDFQD1 \entry_reg[14][3]  ( .D(N10320), .E(N10363), .CP(clk), .Q(
        \entry[14][3] ) );
  EDFQD1 \entry_reg[14][2]  ( .D(N10319), .E(N10363), .CP(clk), .Q(
        \entry[14][2] ) );
  EDFQD1 \entry_reg[14][1]  ( .D(N10318), .E(N10363), .CP(clk), .Q(
        \entry[14][1] ) );
  EDFQD1 \entry_reg[14][0]  ( .D(N10317), .E(N10363), .CP(clk), .Q(
        \entry[14][0] ) );
  EDFQD1 \entry_reg[13][31]  ( .D(N10348), .E(N10362), .CP(clk), .Q(
        \entry[13][31] ) );
  EDFQD1 \entry_reg[13][30]  ( .D(N10347), .E(N10362), .CP(clk), .Q(
        \entry[13][30] ) );
  EDFQD1 \entry_reg[13][29]  ( .D(N10346), .E(N10362), .CP(clk), .Q(
        \entry[13][29] ) );
  EDFQD1 \entry_reg[13][28]  ( .D(N10345), .E(N10362), .CP(clk), .Q(
        \entry[13][28] ) );
  EDFQD1 \entry_reg[13][27]  ( .D(N10344), .E(N10362), .CP(clk), .Q(
        \entry[13][27] ) );
  EDFQD1 \entry_reg[13][26]  ( .D(N10343), .E(N10362), .CP(clk), .Q(
        \entry[13][26] ) );
  EDFQD1 \entry_reg[13][25]  ( .D(N10342), .E(N10362), .CP(clk), .Q(
        \entry[13][25] ) );
  EDFQD1 \entry_reg[13][24]  ( .D(N10341), .E(N10362), .CP(clk), .Q(
        \entry[13][24] ) );
  EDFQD1 \entry_reg[13][23]  ( .D(N10340), .E(N10362), .CP(clk), .Q(
        \entry[13][23] ) );
  EDFQD1 \entry_reg[13][22]  ( .D(N10339), .E(N10362), .CP(clk), .Q(
        \entry[13][22] ) );
  EDFQD1 \entry_reg[13][21]  ( .D(N10338), .E(N10362), .CP(clk), .Q(
        \entry[13][21] ) );
  EDFQD1 \entry_reg[13][20]  ( .D(N10337), .E(N10362), .CP(clk), .Q(
        \entry[13][20] ) );
  EDFQD1 \entry_reg[13][19]  ( .D(N10336), .E(N10362), .CP(clk), .Q(
        \entry[13][19] ) );
  EDFQD1 \entry_reg[13][18]  ( .D(N10335), .E(N10362), .CP(clk), .Q(
        \entry[13][18] ) );
  EDFQD1 \entry_reg[13][17]  ( .D(N10334), .E(N10362), .CP(clk), .Q(
        \entry[13][17] ) );
  EDFQD1 \entry_reg[13][16]  ( .D(N10333), .E(N10362), .CP(clk), .Q(
        \entry[13][16] ) );
  EDFQD1 \entry_reg[13][15]  ( .D(N10332), .E(N10362), .CP(clk), .Q(
        \entry[13][15] ) );
  EDFQD1 \entry_reg[13][14]  ( .D(N10331), .E(N10362), .CP(clk), .Q(
        \entry[13][14] ) );
  EDFQD1 \entry_reg[13][13]  ( .D(N10330), .E(N10362), .CP(clk), .Q(
        \entry[13][13] ) );
  EDFQD1 \entry_reg[13][12]  ( .D(N10329), .E(N10362), .CP(clk), .Q(
        \entry[13][12] ) );
  EDFQD1 \entry_reg[13][11]  ( .D(N10328), .E(N10362), .CP(clk), .Q(
        \entry[13][11] ) );
  EDFQD1 \entry_reg[13][10]  ( .D(N10327), .E(N10362), .CP(clk), .Q(
        \entry[13][10] ) );
  EDFQD1 \entry_reg[13][9]  ( .D(N10326), .E(N10362), .CP(clk), .Q(
        \entry[13][9] ) );
  EDFQD1 \entry_reg[13][8]  ( .D(N10325), .E(N10362), .CP(clk), .Q(
        \entry[13][8] ) );
  EDFQD1 \entry_reg[13][7]  ( .D(N10324), .E(N10362), .CP(clk), .Q(
        \entry[13][7] ) );
  EDFQD1 \entry_reg[13][6]  ( .D(N10323), .E(N10362), .CP(clk), .Q(
        \entry[13][6] ) );
  EDFQD1 \entry_reg[13][5]  ( .D(N10322), .E(N10362), .CP(clk), .Q(
        \entry[13][5] ) );
  EDFQD1 \entry_reg[13][4]  ( .D(N10321), .E(N10362), .CP(clk), .Q(
        \entry[13][4] ) );
  EDFQD1 \entry_reg[13][3]  ( .D(N10320), .E(N10362), .CP(clk), .Q(
        \entry[13][3] ) );
  EDFQD1 \entry_reg[13][2]  ( .D(N10319), .E(N10362), .CP(clk), .Q(
        \entry[13][2] ) );
  EDFQD1 \entry_reg[13][1]  ( .D(N10318), .E(N10362), .CP(clk), .Q(
        \entry[13][1] ) );
  EDFQD1 \entry_reg[13][0]  ( .D(N10317), .E(N10362), .CP(clk), .Q(
        \entry[13][0] ) );
  EDFQD1 \entry_reg[12][31]  ( .D(N10348), .E(N10361), .CP(clk), .Q(
        \entry[12][31] ) );
  EDFQD1 \entry_reg[12][30]  ( .D(N10347), .E(N10361), .CP(clk), .Q(
        \entry[12][30] ) );
  EDFQD1 \entry_reg[12][29]  ( .D(N10346), .E(N10361), .CP(clk), .Q(
        \entry[12][29] ) );
  EDFQD1 \entry_reg[12][28]  ( .D(N10345), .E(N10361), .CP(clk), .Q(
        \entry[12][28] ) );
  EDFQD1 \entry_reg[12][27]  ( .D(N10344), .E(N10361), .CP(clk), .Q(
        \entry[12][27] ) );
  EDFQD1 \entry_reg[12][26]  ( .D(N10343), .E(N10361), .CP(clk), .Q(
        \entry[12][26] ) );
  EDFQD1 \entry_reg[12][25]  ( .D(N10342), .E(N10361), .CP(clk), .Q(
        \entry[12][25] ) );
  EDFQD1 \entry_reg[12][24]  ( .D(N10341), .E(N10361), .CP(clk), .Q(
        \entry[12][24] ) );
  EDFQD1 \entry_reg[12][23]  ( .D(N10340), .E(N10361), .CP(clk), .Q(
        \entry[12][23] ) );
  EDFQD1 \entry_reg[12][22]  ( .D(N10339), .E(N10361), .CP(clk), .Q(
        \entry[12][22] ) );
  EDFQD1 \entry_reg[12][21]  ( .D(N10338), .E(N10361), .CP(clk), .Q(
        \entry[12][21] ) );
  EDFQD1 \entry_reg[12][20]  ( .D(N10337), .E(N10361), .CP(clk), .Q(
        \entry[12][20] ) );
  EDFQD1 \entry_reg[12][19]  ( .D(N10336), .E(N10361), .CP(clk), .Q(
        \entry[12][19] ) );
  EDFQD1 \entry_reg[12][18]  ( .D(N10335), .E(N10361), .CP(clk), .Q(
        \entry[12][18] ) );
  EDFQD1 \entry_reg[12][17]  ( .D(N10334), .E(N10361), .CP(clk), .Q(
        \entry[12][17] ) );
  EDFQD1 \entry_reg[12][16]  ( .D(N10333), .E(N10361), .CP(clk), .Q(
        \entry[12][16] ) );
  EDFQD1 \entry_reg[12][15]  ( .D(N10332), .E(N10361), .CP(clk), .Q(
        \entry[12][15] ) );
  EDFQD1 \entry_reg[12][14]  ( .D(N10331), .E(N10361), .CP(clk), .Q(
        \entry[12][14] ) );
  EDFQD1 \entry_reg[12][13]  ( .D(N10330), .E(N10361), .CP(clk), .Q(
        \entry[12][13] ) );
  EDFQD1 \entry_reg[12][12]  ( .D(N10329), .E(N10361), .CP(clk), .Q(
        \entry[12][12] ) );
  EDFQD1 \entry_reg[12][11]  ( .D(N10328), .E(N10361), .CP(clk), .Q(
        \entry[12][11] ) );
  EDFQD1 \entry_reg[12][10]  ( .D(N10327), .E(N10361), .CP(clk), .Q(
        \entry[12][10] ) );
  EDFQD1 \entry_reg[12][9]  ( .D(N10326), .E(N10361), .CP(clk), .Q(
        \entry[12][9] ) );
  EDFQD1 \entry_reg[12][8]  ( .D(N10325), .E(N10361), .CP(clk), .Q(
        \entry[12][8] ) );
  EDFQD1 \entry_reg[12][7]  ( .D(N10324), .E(N10361), .CP(clk), .Q(
        \entry[12][7] ) );
  EDFQD1 \entry_reg[12][6]  ( .D(N10323), .E(N10361), .CP(clk), .Q(
        \entry[12][6] ) );
  EDFQD1 \entry_reg[12][5]  ( .D(N10322), .E(N10361), .CP(clk), .Q(
        \entry[12][5] ) );
  EDFQD1 \entry_reg[12][4]  ( .D(N10321), .E(N10361), .CP(clk), .Q(
        \entry[12][4] ) );
  EDFQD1 \entry_reg[12][3]  ( .D(N10320), .E(N10361), .CP(clk), .Q(
        \entry[12][3] ) );
  EDFQD1 \entry_reg[12][2]  ( .D(N10319), .E(N10361), .CP(clk), .Q(
        \entry[12][2] ) );
  EDFQD1 \entry_reg[12][1]  ( .D(N10318), .E(N10361), .CP(clk), .Q(
        \entry[12][1] ) );
  EDFQD1 \entry_reg[12][0]  ( .D(N10317), .E(N10361), .CP(clk), .Q(
        \entry[12][0] ) );
  EDFQD1 \entry_reg[11][31]  ( .D(N10348), .E(N10360), .CP(clk), .Q(
        \entry[11][31] ) );
  EDFQD1 \entry_reg[11][30]  ( .D(N10347), .E(N10360), .CP(clk), .Q(
        \entry[11][30] ) );
  EDFQD1 \entry_reg[11][29]  ( .D(N10346), .E(N10360), .CP(clk), .Q(
        \entry[11][29] ) );
  EDFQD1 \entry_reg[11][28]  ( .D(N10345), .E(N10360), .CP(clk), .Q(
        \entry[11][28] ) );
  EDFQD1 \entry_reg[11][27]  ( .D(N10344), .E(N10360), .CP(clk), .Q(
        \entry[11][27] ) );
  EDFQD1 \entry_reg[11][26]  ( .D(N10343), .E(N10360), .CP(clk), .Q(
        \entry[11][26] ) );
  EDFQD1 \entry_reg[11][25]  ( .D(N10342), .E(N10360), .CP(clk), .Q(
        \entry[11][25] ) );
  EDFQD1 \entry_reg[11][24]  ( .D(N10341), .E(N10360), .CP(clk), .Q(
        \entry[11][24] ) );
  EDFQD1 \entry_reg[11][23]  ( .D(N10340), .E(N10360), .CP(clk), .Q(
        \entry[11][23] ) );
  EDFQD1 \entry_reg[11][22]  ( .D(N10339), .E(N10360), .CP(clk), .Q(
        \entry[11][22] ) );
  EDFQD1 \entry_reg[11][21]  ( .D(N10338), .E(N10360), .CP(clk), .Q(
        \entry[11][21] ) );
  EDFQD1 \entry_reg[11][20]  ( .D(N10337), .E(N10360), .CP(clk), .Q(
        \entry[11][20] ) );
  EDFQD1 \entry_reg[11][19]  ( .D(N10336), .E(N10360), .CP(clk), .Q(
        \entry[11][19] ) );
  EDFQD1 \entry_reg[11][18]  ( .D(N10335), .E(N10360), .CP(clk), .Q(
        \entry[11][18] ) );
  EDFQD1 \entry_reg[11][17]  ( .D(N10334), .E(N10360), .CP(clk), .Q(
        \entry[11][17] ) );
  EDFQD1 \entry_reg[11][16]  ( .D(N10333), .E(N10360), .CP(clk), .Q(
        \entry[11][16] ) );
  EDFQD1 \entry_reg[11][15]  ( .D(N10332), .E(N10360), .CP(clk), .Q(
        \entry[11][15] ) );
  EDFQD1 \entry_reg[11][14]  ( .D(N10331), .E(N10360), .CP(clk), .Q(
        \entry[11][14] ) );
  EDFQD1 \entry_reg[11][13]  ( .D(N10330), .E(N10360), .CP(clk), .Q(
        \entry[11][13] ) );
  EDFQD1 \entry_reg[11][12]  ( .D(N10329), .E(N10360), .CP(clk), .Q(
        \entry[11][12] ) );
  EDFQD1 \entry_reg[11][11]  ( .D(N10328), .E(N10360), .CP(clk), .Q(
        \entry[11][11] ) );
  EDFQD1 \entry_reg[11][10]  ( .D(N10327), .E(N10360), .CP(clk), .Q(
        \entry[11][10] ) );
  EDFQD1 \entry_reg[11][9]  ( .D(N10326), .E(N10360), .CP(clk), .Q(
        \entry[11][9] ) );
  EDFQD1 \entry_reg[11][8]  ( .D(N10325), .E(N10360), .CP(clk), .Q(
        \entry[11][8] ) );
  EDFQD1 \entry_reg[11][7]  ( .D(N10324), .E(N10360), .CP(clk), .Q(
        \entry[11][7] ) );
  EDFQD1 \entry_reg[11][6]  ( .D(N10323), .E(N10360), .CP(clk), .Q(
        \entry[11][6] ) );
  EDFQD1 \entry_reg[11][5]  ( .D(N10322), .E(N10360), .CP(clk), .Q(
        \entry[11][5] ) );
  EDFQD1 \entry_reg[11][4]  ( .D(N10321), .E(N10360), .CP(clk), .Q(
        \entry[11][4] ) );
  EDFQD1 \entry_reg[11][3]  ( .D(N10320), .E(N10360), .CP(clk), .Q(
        \entry[11][3] ) );
  EDFQD1 \entry_reg[11][2]  ( .D(N10319), .E(N10360), .CP(clk), .Q(
        \entry[11][2] ) );
  EDFQD1 \entry_reg[11][1]  ( .D(N10318), .E(N10360), .CP(clk), .Q(
        \entry[11][1] ) );
  EDFQD1 \entry_reg[11][0]  ( .D(N10317), .E(N10360), .CP(clk), .Q(
        \entry[11][0] ) );
  EDFQD1 \entry_reg[10][31]  ( .D(N10348), .E(N10359), .CP(clk), .Q(
        \entry[10][31] ) );
  EDFQD1 \entry_reg[10][30]  ( .D(N10347), .E(N10359), .CP(clk), .Q(
        \entry[10][30] ) );
  EDFQD1 \entry_reg[10][29]  ( .D(N10346), .E(N10359), .CP(clk), .Q(
        \entry[10][29] ) );
  EDFQD1 \entry_reg[10][28]  ( .D(N10345), .E(N10359), .CP(clk), .Q(
        \entry[10][28] ) );
  EDFQD1 \entry_reg[10][27]  ( .D(N10344), .E(N10359), .CP(clk), .Q(
        \entry[10][27] ) );
  EDFQD1 \entry_reg[10][26]  ( .D(N10343), .E(N10359), .CP(clk), .Q(
        \entry[10][26] ) );
  EDFQD1 \entry_reg[10][25]  ( .D(N10342), .E(N10359), .CP(clk), .Q(
        \entry[10][25] ) );
  EDFQD1 \entry_reg[10][24]  ( .D(N10341), .E(N10359), .CP(clk), .Q(
        \entry[10][24] ) );
  EDFQD1 \entry_reg[10][23]  ( .D(N10340), .E(N10359), .CP(clk), .Q(
        \entry[10][23] ) );
  EDFQD1 \entry_reg[10][22]  ( .D(N10339), .E(N10359), .CP(clk), .Q(
        \entry[10][22] ) );
  EDFQD1 \entry_reg[10][21]  ( .D(N10338), .E(N10359), .CP(clk), .Q(
        \entry[10][21] ) );
  EDFQD1 \entry_reg[10][20]  ( .D(N10337), .E(N10359), .CP(clk), .Q(
        \entry[10][20] ) );
  EDFQD1 \entry_reg[10][19]  ( .D(N10336), .E(N10359), .CP(clk), .Q(
        \entry[10][19] ) );
  EDFQD1 \entry_reg[10][18]  ( .D(N10335), .E(N10359), .CP(clk), .Q(
        \entry[10][18] ) );
  EDFQD1 \entry_reg[10][17]  ( .D(N10334), .E(N10359), .CP(clk), .Q(
        \entry[10][17] ) );
  EDFQD1 \entry_reg[10][16]  ( .D(N10333), .E(N10359), .CP(clk), .Q(
        \entry[10][16] ) );
  EDFQD1 \entry_reg[10][15]  ( .D(N10332), .E(N10359), .CP(clk), .Q(
        \entry[10][15] ) );
  EDFQD1 \entry_reg[10][14]  ( .D(N10331), .E(N10359), .CP(clk), .Q(
        \entry[10][14] ) );
  EDFQD1 \entry_reg[10][13]  ( .D(N10330), .E(N10359), .CP(clk), .Q(
        \entry[10][13] ) );
  EDFQD1 \entry_reg[10][12]  ( .D(N10329), .E(N10359), .CP(clk), .Q(
        \entry[10][12] ) );
  EDFQD1 \entry_reg[10][11]  ( .D(N10328), .E(N10359), .CP(clk), .Q(
        \entry[10][11] ) );
  EDFQD1 \entry_reg[10][10]  ( .D(N10327), .E(N10359), .CP(clk), .Q(
        \entry[10][10] ) );
  EDFQD1 \entry_reg[10][9]  ( .D(N10326), .E(N10359), .CP(clk), .Q(
        \entry[10][9] ) );
  EDFQD1 \entry_reg[10][8]  ( .D(N10325), .E(N10359), .CP(clk), .Q(
        \entry[10][8] ) );
  EDFQD1 \entry_reg[10][7]  ( .D(N10324), .E(N10359), .CP(clk), .Q(
        \entry[10][7] ) );
  EDFQD1 \entry_reg[10][6]  ( .D(N10323), .E(N10359), .CP(clk), .Q(
        \entry[10][6] ) );
  EDFQD1 \entry_reg[10][5]  ( .D(N10322), .E(N10359), .CP(clk), .Q(
        \entry[10][5] ) );
  EDFQD1 \entry_reg[10][4]  ( .D(N10321), .E(N10359), .CP(clk), .Q(
        \entry[10][4] ) );
  EDFQD1 \entry_reg[10][3]  ( .D(N10320), .E(N10359), .CP(clk), .Q(
        \entry[10][3] ) );
  EDFQD1 \entry_reg[10][2]  ( .D(N10319), .E(N10359), .CP(clk), .Q(
        \entry[10][2] ) );
  EDFQD1 \entry_reg[10][1]  ( .D(N10318), .E(N10359), .CP(clk), .Q(
        \entry[10][1] ) );
  EDFQD1 \entry_reg[10][0]  ( .D(N10317), .E(N10359), .CP(clk), .Q(
        \entry[10][0] ) );
  EDFQD1 \entry_reg[9][31]  ( .D(N10348), .E(N10358), .CP(clk), .Q(
        \entry[9][31] ) );
  EDFQD1 \entry_reg[9][30]  ( .D(N10347), .E(N10358), .CP(clk), .Q(
        \entry[9][30] ) );
  EDFQD1 \entry_reg[9][29]  ( .D(N10346), .E(N10358), .CP(clk), .Q(
        \entry[9][29] ) );
  EDFQD1 \entry_reg[9][28]  ( .D(N10345), .E(N10358), .CP(clk), .Q(
        \entry[9][28] ) );
  EDFQD1 \entry_reg[9][27]  ( .D(N10344), .E(N10358), .CP(clk), .Q(
        \entry[9][27] ) );
  EDFQD1 \entry_reg[9][26]  ( .D(N10343), .E(N10358), .CP(clk), .Q(
        \entry[9][26] ) );
  EDFQD1 \entry_reg[9][25]  ( .D(N10342), .E(N10358), .CP(clk), .Q(
        \entry[9][25] ) );
  EDFQD1 \entry_reg[9][24]  ( .D(N10341), .E(N10358), .CP(clk), .Q(
        \entry[9][24] ) );
  EDFQD1 \entry_reg[9][23]  ( .D(N10340), .E(N10358), .CP(clk), .Q(
        \entry[9][23] ) );
  EDFQD1 \entry_reg[9][22]  ( .D(N10339), .E(N10358), .CP(clk), .Q(
        \entry[9][22] ) );
  EDFQD1 \entry_reg[9][21]  ( .D(N10338), .E(N10358), .CP(clk), .Q(
        \entry[9][21] ) );
  EDFQD1 \entry_reg[9][20]  ( .D(N10337), .E(N10358), .CP(clk), .Q(
        \entry[9][20] ) );
  EDFQD1 \entry_reg[9][19]  ( .D(N10336), .E(N10358), .CP(clk), .Q(
        \entry[9][19] ) );
  EDFQD1 \entry_reg[9][18]  ( .D(N10335), .E(N10358), .CP(clk), .Q(
        \entry[9][18] ) );
  EDFQD1 \entry_reg[9][17]  ( .D(N10334), .E(N10358), .CP(clk), .Q(
        \entry[9][17] ) );
  EDFQD1 \entry_reg[9][16]  ( .D(N10333), .E(N10358), .CP(clk), .Q(
        \entry[9][16] ) );
  EDFQD1 \entry_reg[9][15]  ( .D(N10332), .E(N10358), .CP(clk), .Q(
        \entry[9][15] ) );
  EDFQD1 \entry_reg[9][14]  ( .D(N10331), .E(N10358), .CP(clk), .Q(
        \entry[9][14] ) );
  EDFQD1 \entry_reg[9][13]  ( .D(N10330), .E(N10358), .CP(clk), .Q(
        \entry[9][13] ) );
  EDFQD1 \entry_reg[9][12]  ( .D(N10329), .E(N10358), .CP(clk), .Q(
        \entry[9][12] ) );
  EDFQD1 \entry_reg[9][11]  ( .D(N10328), .E(N10358), .CP(clk), .Q(
        \entry[9][11] ) );
  EDFQD1 \entry_reg[9][10]  ( .D(N10327), .E(N10358), .CP(clk), .Q(
        \entry[9][10] ) );
  EDFQD1 \entry_reg[9][9]  ( .D(N10326), .E(N10358), .CP(clk), .Q(
        \entry[9][9] ) );
  EDFQD1 \entry_reg[9][8]  ( .D(N10325), .E(N10358), .CP(clk), .Q(
        \entry[9][8] ) );
  EDFQD1 \entry_reg[9][7]  ( .D(N10324), .E(N10358), .CP(clk), .Q(
        \entry[9][7] ) );
  EDFQD1 \entry_reg[9][6]  ( .D(N10323), .E(N10358), .CP(clk), .Q(
        \entry[9][6] ) );
  EDFQD1 \entry_reg[9][5]  ( .D(N10322), .E(N10358), .CP(clk), .Q(
        \entry[9][5] ) );
  EDFQD1 \entry_reg[9][4]  ( .D(N10321), .E(N10358), .CP(clk), .Q(
        \entry[9][4] ) );
  EDFQD1 \entry_reg[9][3]  ( .D(N10320), .E(N10358), .CP(clk), .Q(
        \entry[9][3] ) );
  EDFQD1 \entry_reg[9][2]  ( .D(N10319), .E(N10358), .CP(clk), .Q(
        \entry[9][2] ) );
  EDFQD1 \entry_reg[9][1]  ( .D(N10318), .E(N10358), .CP(clk), .Q(
        \entry[9][1] ) );
  EDFQD1 \entry_reg[9][0]  ( .D(N10317), .E(N10358), .CP(clk), .Q(
        \entry[9][0] ) );
  EDFQD1 \entry_reg[8][31]  ( .D(N10348), .E(N10357), .CP(clk), .Q(
        \entry[8][31] ) );
  EDFQD1 \entry_reg[8][30]  ( .D(N10347), .E(N10357), .CP(clk), .Q(
        \entry[8][30] ) );
  EDFQD1 \entry_reg[8][29]  ( .D(N10346), .E(N10357), .CP(clk), .Q(
        \entry[8][29] ) );
  EDFQD1 \entry_reg[8][28]  ( .D(N10345), .E(N10357), .CP(clk), .Q(
        \entry[8][28] ) );
  EDFQD1 \entry_reg[8][27]  ( .D(N10344), .E(N10357), .CP(clk), .Q(
        \entry[8][27] ) );
  EDFQD1 \entry_reg[8][26]  ( .D(N10343), .E(N10357), .CP(clk), .Q(
        \entry[8][26] ) );
  EDFQD1 \entry_reg[8][25]  ( .D(N10342), .E(N10357), .CP(clk), .Q(
        \entry[8][25] ) );
  EDFQD1 \entry_reg[8][24]  ( .D(N10341), .E(N10357), .CP(clk), .Q(
        \entry[8][24] ) );
  EDFQD1 \entry_reg[8][23]  ( .D(N10340), .E(N10357), .CP(clk), .Q(
        \entry[8][23] ) );
  EDFQD1 \entry_reg[8][22]  ( .D(N10339), .E(N10357), .CP(clk), .Q(
        \entry[8][22] ) );
  EDFQD1 \entry_reg[8][21]  ( .D(N10338), .E(N10357), .CP(clk), .Q(
        \entry[8][21] ) );
  EDFQD1 \entry_reg[8][20]  ( .D(N10337), .E(N10357), .CP(clk), .Q(
        \entry[8][20] ) );
  EDFQD1 \entry_reg[8][19]  ( .D(N10336), .E(N10357), .CP(clk), .Q(
        \entry[8][19] ) );
  EDFQD1 \entry_reg[8][18]  ( .D(N10335), .E(N10357), .CP(clk), .Q(
        \entry[8][18] ) );
  EDFQD1 \entry_reg[8][17]  ( .D(N10334), .E(N10357), .CP(clk), .Q(
        \entry[8][17] ) );
  EDFQD1 \entry_reg[8][16]  ( .D(N10333), .E(N10357), .CP(clk), .Q(
        \entry[8][16] ) );
  EDFQD1 \entry_reg[8][15]  ( .D(N10332), .E(N10357), .CP(clk), .Q(
        \entry[8][15] ) );
  EDFQD1 \entry_reg[8][14]  ( .D(N10331), .E(N10357), .CP(clk), .Q(
        \entry[8][14] ) );
  EDFQD1 \entry_reg[8][13]  ( .D(N10330), .E(N10357), .CP(clk), .Q(
        \entry[8][13] ) );
  EDFQD1 \entry_reg[8][12]  ( .D(N10329), .E(N10357), .CP(clk), .Q(
        \entry[8][12] ) );
  EDFQD1 \entry_reg[8][11]  ( .D(N10328), .E(N10357), .CP(clk), .Q(
        \entry[8][11] ) );
  EDFQD1 \entry_reg[8][10]  ( .D(N10327), .E(N10357), .CP(clk), .Q(
        \entry[8][10] ) );
  EDFQD1 \entry_reg[8][9]  ( .D(N10326), .E(N10357), .CP(clk), .Q(
        \entry[8][9] ) );
  EDFQD1 \entry_reg[8][8]  ( .D(N10325), .E(N10357), .CP(clk), .Q(
        \entry[8][8] ) );
  EDFQD1 \entry_reg[8][7]  ( .D(N10324), .E(N10357), .CP(clk), .Q(
        \entry[8][7] ) );
  EDFQD1 \entry_reg[8][6]  ( .D(N10323), .E(N10357), .CP(clk), .Q(
        \entry[8][6] ) );
  EDFQD1 \entry_reg[8][5]  ( .D(N10322), .E(N10357), .CP(clk), .Q(
        \entry[8][5] ) );
  EDFQD1 \entry_reg[8][4]  ( .D(N10321), .E(N10357), .CP(clk), .Q(
        \entry[8][4] ) );
  EDFQD1 \entry_reg[8][3]  ( .D(N10320), .E(N10357), .CP(clk), .Q(
        \entry[8][3] ) );
  EDFQD1 \entry_reg[8][2]  ( .D(N10319), .E(N10357), .CP(clk), .Q(
        \entry[8][2] ) );
  EDFQD1 \entry_reg[8][1]  ( .D(N10318), .E(N10357), .CP(clk), .Q(
        \entry[8][1] ) );
  EDFQD1 \entry_reg[8][0]  ( .D(N10317), .E(N10357), .CP(clk), .Q(
        \entry[8][0] ) );
  EDFQD1 \entry_reg[7][31]  ( .D(N10348), .E(N10356), .CP(clk), .Q(
        \entry[7][31] ) );
  EDFQD1 \entry_reg[7][30]  ( .D(N10347), .E(N10356), .CP(clk), .Q(
        \entry[7][30] ) );
  EDFQD1 \entry_reg[7][29]  ( .D(N10346), .E(N10356), .CP(clk), .Q(
        \entry[7][29] ) );
  EDFQD1 \entry_reg[7][28]  ( .D(N10345), .E(N10356), .CP(clk), .Q(
        \entry[7][28] ) );
  EDFQD1 \entry_reg[7][27]  ( .D(N10344), .E(N10356), .CP(clk), .Q(
        \entry[7][27] ) );
  EDFQD1 \entry_reg[7][26]  ( .D(N10343), .E(N10356), .CP(clk), .Q(
        \entry[7][26] ) );
  EDFQD1 \entry_reg[7][25]  ( .D(N10342), .E(N10356), .CP(clk), .Q(
        \entry[7][25] ) );
  EDFQD1 \entry_reg[7][24]  ( .D(N10341), .E(N10356), .CP(clk), .Q(
        \entry[7][24] ) );
  EDFQD1 \entry_reg[7][23]  ( .D(N10340), .E(N10356), .CP(clk), .Q(
        \entry[7][23] ) );
  EDFQD1 \entry_reg[7][22]  ( .D(N10339), .E(N10356), .CP(clk), .Q(
        \entry[7][22] ) );
  EDFQD1 \entry_reg[7][21]  ( .D(N10338), .E(N10356), .CP(clk), .Q(
        \entry[7][21] ) );
  EDFQD1 \entry_reg[7][20]  ( .D(N10337), .E(N10356), .CP(clk), .Q(
        \entry[7][20] ) );
  EDFQD1 \entry_reg[7][19]  ( .D(N10336), .E(N10356), .CP(clk), .Q(
        \entry[7][19] ) );
  EDFQD1 \entry_reg[7][18]  ( .D(N10335), .E(N10356), .CP(clk), .Q(
        \entry[7][18] ) );
  EDFQD1 \entry_reg[7][17]  ( .D(N10334), .E(N10356), .CP(clk), .Q(
        \entry[7][17] ) );
  EDFQD1 \entry_reg[7][16]  ( .D(N10333), .E(N10356), .CP(clk), .Q(
        \entry[7][16] ) );
  EDFQD1 \entry_reg[7][15]  ( .D(N10332), .E(N10356), .CP(clk), .Q(
        \entry[7][15] ) );
  EDFQD1 \entry_reg[7][14]  ( .D(N10331), .E(N10356), .CP(clk), .Q(
        \entry[7][14] ) );
  EDFQD1 \entry_reg[7][13]  ( .D(N10330), .E(N10356), .CP(clk), .Q(
        \entry[7][13] ) );
  EDFQD1 \entry_reg[7][12]  ( .D(N10329), .E(N10356), .CP(clk), .Q(
        \entry[7][12] ) );
  EDFQD1 \entry_reg[7][11]  ( .D(N10328), .E(N10356), .CP(clk), .Q(
        \entry[7][11] ) );
  EDFQD1 \entry_reg[7][10]  ( .D(N10327), .E(N10356), .CP(clk), .Q(
        \entry[7][10] ) );
  EDFQD1 \entry_reg[7][9]  ( .D(N10326), .E(N10356), .CP(clk), .Q(
        \entry[7][9] ) );
  EDFQD1 \entry_reg[7][8]  ( .D(N10325), .E(N10356), .CP(clk), .Q(
        \entry[7][8] ) );
  EDFQD1 \entry_reg[7][7]  ( .D(N10324), .E(N10356), .CP(clk), .Q(
        \entry[7][7] ) );
  EDFQD1 \entry_reg[7][6]  ( .D(N10323), .E(N10356), .CP(clk), .Q(
        \entry[7][6] ) );
  EDFQD1 \entry_reg[7][5]  ( .D(N10322), .E(N10356), .CP(clk), .Q(
        \entry[7][5] ) );
  EDFQD1 \entry_reg[7][4]  ( .D(N10321), .E(N10356), .CP(clk), .Q(
        \entry[7][4] ) );
  EDFQD1 \entry_reg[7][3]  ( .D(N10320), .E(N10356), .CP(clk), .Q(
        \entry[7][3] ) );
  EDFQD1 \entry_reg[7][2]  ( .D(N10319), .E(N10356), .CP(clk), .Q(
        \entry[7][2] ) );
  EDFQD1 \entry_reg[7][1]  ( .D(N10318), .E(N10356), .CP(clk), .Q(
        \entry[7][1] ) );
  EDFQD1 \entry_reg[7][0]  ( .D(N10317), .E(N10356), .CP(clk), .Q(
        \entry[7][0] ) );
  EDFQD1 \entry_reg[6][31]  ( .D(N10348), .E(N10355), .CP(clk), .Q(
        \entry[6][31] ) );
  EDFQD1 \entry_reg[6][30]  ( .D(N10347), .E(N10355), .CP(clk), .Q(
        \entry[6][30] ) );
  EDFQD1 \entry_reg[6][29]  ( .D(N10346), .E(N10355), .CP(clk), .Q(
        \entry[6][29] ) );
  EDFQD1 \entry_reg[6][28]  ( .D(N10345), .E(N10355), .CP(clk), .Q(
        \entry[6][28] ) );
  EDFQD1 \entry_reg[6][27]  ( .D(N10344), .E(N10355), .CP(clk), .Q(
        \entry[6][27] ) );
  EDFQD1 \entry_reg[6][26]  ( .D(N10343), .E(N10355), .CP(clk), .Q(
        \entry[6][26] ) );
  EDFQD1 \entry_reg[6][25]  ( .D(N10342), .E(N10355), .CP(clk), .Q(
        \entry[6][25] ) );
  EDFQD1 \entry_reg[6][24]  ( .D(N10341), .E(N10355), .CP(clk), .Q(
        \entry[6][24] ) );
  EDFQD1 \entry_reg[6][23]  ( .D(N10340), .E(N10355), .CP(clk), .Q(
        \entry[6][23] ) );
  EDFQD1 \entry_reg[6][22]  ( .D(N10339), .E(N10355), .CP(clk), .Q(
        \entry[6][22] ) );
  EDFQD1 \entry_reg[6][21]  ( .D(N10338), .E(N10355), .CP(clk), .Q(
        \entry[6][21] ) );
  EDFQD1 \entry_reg[6][20]  ( .D(N10337), .E(N10355), .CP(clk), .Q(
        \entry[6][20] ) );
  EDFQD1 \entry_reg[6][19]  ( .D(N10336), .E(N10355), .CP(clk), .Q(
        \entry[6][19] ) );
  EDFQD1 \entry_reg[6][18]  ( .D(N10335), .E(N10355), .CP(clk), .Q(
        \entry[6][18] ) );
  EDFQD1 \entry_reg[6][17]  ( .D(N10334), .E(N10355), .CP(clk), .Q(
        \entry[6][17] ) );
  EDFQD1 \entry_reg[6][16]  ( .D(N10333), .E(N10355), .CP(clk), .Q(
        \entry[6][16] ) );
  EDFQD1 \entry_reg[6][15]  ( .D(N10332), .E(N10355), .CP(clk), .Q(
        \entry[6][15] ) );
  EDFQD1 \entry_reg[6][14]  ( .D(N10331), .E(N10355), .CP(clk), .Q(
        \entry[6][14] ) );
  EDFQD1 \entry_reg[6][13]  ( .D(N10330), .E(N10355), .CP(clk), .Q(
        \entry[6][13] ) );
  EDFQD1 \entry_reg[6][12]  ( .D(N10329), .E(N10355), .CP(clk), .Q(
        \entry[6][12] ) );
  EDFQD1 \entry_reg[6][11]  ( .D(N10328), .E(N10355), .CP(clk), .Q(
        \entry[6][11] ) );
  EDFQD1 \entry_reg[6][10]  ( .D(N10327), .E(N10355), .CP(clk), .Q(
        \entry[6][10] ) );
  EDFQD1 \entry_reg[6][9]  ( .D(N10326), .E(N10355), .CP(clk), .Q(
        \entry[6][9] ) );
  EDFQD1 \entry_reg[6][8]  ( .D(N10325), .E(N10355), .CP(clk), .Q(
        \entry[6][8] ) );
  EDFQD1 \entry_reg[6][7]  ( .D(N10324), .E(N10355), .CP(clk), .Q(
        \entry[6][7] ) );
  EDFQD1 \entry_reg[6][6]  ( .D(N10323), .E(N10355), .CP(clk), .Q(
        \entry[6][6] ) );
  EDFQD1 \entry_reg[6][5]  ( .D(N10322), .E(N10355), .CP(clk), .Q(
        \entry[6][5] ) );
  EDFQD1 \entry_reg[6][4]  ( .D(N10321), .E(N10355), .CP(clk), .Q(
        \entry[6][4] ) );
  EDFQD1 \entry_reg[6][3]  ( .D(N10320), .E(N10355), .CP(clk), .Q(
        \entry[6][3] ) );
  EDFQD1 \entry_reg[6][2]  ( .D(N10319), .E(N10355), .CP(clk), .Q(
        \entry[6][2] ) );
  EDFQD1 \entry_reg[6][1]  ( .D(N10318), .E(N10355), .CP(clk), .Q(
        \entry[6][1] ) );
  EDFQD1 \entry_reg[6][0]  ( .D(N10317), .E(N10355), .CP(clk), .Q(
        \entry[6][0] ) );
  EDFQD1 \entry_reg[5][31]  ( .D(N10348), .E(N10354), .CP(clk), .Q(
        \entry[5][31] ) );
  EDFQD1 \entry_reg[5][30]  ( .D(N10347), .E(N10354), .CP(clk), .Q(
        \entry[5][30] ) );
  EDFQD1 \entry_reg[5][29]  ( .D(N10346), .E(N10354), .CP(clk), .Q(
        \entry[5][29] ) );
  EDFQD1 \entry_reg[5][28]  ( .D(N10345), .E(N10354), .CP(clk), .Q(
        \entry[5][28] ) );
  EDFQD1 \entry_reg[5][27]  ( .D(N10344), .E(N10354), .CP(clk), .Q(
        \entry[5][27] ) );
  EDFQD1 \entry_reg[5][26]  ( .D(N10343), .E(N10354), .CP(clk), .Q(
        \entry[5][26] ) );
  EDFQD1 \entry_reg[5][25]  ( .D(N10342), .E(N10354), .CP(clk), .Q(
        \entry[5][25] ) );
  EDFQD1 \entry_reg[5][24]  ( .D(N10341), .E(N10354), .CP(clk), .Q(
        \entry[5][24] ) );
  EDFQD1 \entry_reg[5][23]  ( .D(N10340), .E(N10354), .CP(clk), .Q(
        \entry[5][23] ) );
  EDFQD1 \entry_reg[5][22]  ( .D(N10339), .E(N10354), .CP(clk), .Q(
        \entry[5][22] ) );
  EDFQD1 \entry_reg[5][21]  ( .D(N10338), .E(N10354), .CP(clk), .Q(
        \entry[5][21] ) );
  EDFQD1 \entry_reg[5][20]  ( .D(N10337), .E(N10354), .CP(clk), .Q(
        \entry[5][20] ) );
  EDFQD1 \entry_reg[5][19]  ( .D(N10336), .E(N10354), .CP(clk), .Q(
        \entry[5][19] ) );
  EDFQD1 \entry_reg[5][18]  ( .D(N10335), .E(N10354), .CP(clk), .Q(
        \entry[5][18] ) );
  EDFQD1 \entry_reg[5][17]  ( .D(N10334), .E(N10354), .CP(clk), .Q(
        \entry[5][17] ) );
  EDFQD1 \entry_reg[5][16]  ( .D(N10333), .E(N10354), .CP(clk), .Q(
        \entry[5][16] ) );
  EDFQD1 \entry_reg[5][15]  ( .D(N10332), .E(N10354), .CP(clk), .Q(
        \entry[5][15] ) );
  EDFQD1 \entry_reg[5][14]  ( .D(N10331), .E(N10354), .CP(clk), .Q(
        \entry[5][14] ) );
  EDFQD1 \entry_reg[5][13]  ( .D(N10330), .E(N10354), .CP(clk), .Q(
        \entry[5][13] ) );
  EDFQD1 \entry_reg[5][12]  ( .D(N10329), .E(N10354), .CP(clk), .Q(
        \entry[5][12] ) );
  EDFQD1 \entry_reg[5][11]  ( .D(N10328), .E(N10354), .CP(clk), .Q(
        \entry[5][11] ) );
  EDFQD1 \entry_reg[5][10]  ( .D(N10327), .E(N10354), .CP(clk), .Q(
        \entry[5][10] ) );
  EDFQD1 \entry_reg[5][9]  ( .D(N10326), .E(N10354), .CP(clk), .Q(
        \entry[5][9] ) );
  EDFQD1 \entry_reg[5][8]  ( .D(N10325), .E(N10354), .CP(clk), .Q(
        \entry[5][8] ) );
  EDFQD1 \entry_reg[5][7]  ( .D(N10324), .E(N10354), .CP(clk), .Q(
        \entry[5][7] ) );
  EDFQD1 \entry_reg[5][6]  ( .D(N10323), .E(N10354), .CP(clk), .Q(
        \entry[5][6] ) );
  EDFQD1 \entry_reg[5][5]  ( .D(N10322), .E(N10354), .CP(clk), .Q(
        \entry[5][5] ) );
  EDFQD1 \entry_reg[5][4]  ( .D(N10321), .E(N10354), .CP(clk), .Q(
        \entry[5][4] ) );
  EDFQD1 \entry_reg[5][3]  ( .D(N10320), .E(N10354), .CP(clk), .Q(
        \entry[5][3] ) );
  EDFQD1 \entry_reg[5][2]  ( .D(N10319), .E(N10354), .CP(clk), .Q(
        \entry[5][2] ) );
  EDFQD1 \entry_reg[5][1]  ( .D(N10318), .E(N10354), .CP(clk), .Q(
        \entry[5][1] ) );
  EDFQD1 \entry_reg[5][0]  ( .D(N10317), .E(N10354), .CP(clk), .Q(
        \entry[5][0] ) );
  EDFQD1 \entry_reg[4][31]  ( .D(N10348), .E(N10353), .CP(clk), .Q(
        \entry[4][31] ) );
  EDFQD1 \entry_reg[4][30]  ( .D(N10347), .E(N10353), .CP(clk), .Q(
        \entry[4][30] ) );
  EDFQD1 \entry_reg[4][29]  ( .D(N10346), .E(N10353), .CP(clk), .Q(
        \entry[4][29] ) );
  EDFQD1 \entry_reg[4][28]  ( .D(N10345), .E(N10353), .CP(clk), .Q(
        \entry[4][28] ) );
  EDFQD1 \entry_reg[4][27]  ( .D(N10344), .E(N10353), .CP(clk), .Q(
        \entry[4][27] ) );
  EDFQD1 \entry_reg[4][26]  ( .D(N10343), .E(N10353), .CP(clk), .Q(
        \entry[4][26] ) );
  EDFQD1 \entry_reg[4][25]  ( .D(N10342), .E(N10353), .CP(clk), .Q(
        \entry[4][25] ) );
  EDFQD1 \entry_reg[4][24]  ( .D(N10341), .E(N10353), .CP(clk), .Q(
        \entry[4][24] ) );
  EDFQD1 \entry_reg[4][23]  ( .D(N10340), .E(N10353), .CP(clk), .Q(
        \entry[4][23] ) );
  EDFQD1 \entry_reg[4][22]  ( .D(N10339), .E(N10353), .CP(clk), .Q(
        \entry[4][22] ) );
  EDFQD1 \entry_reg[4][21]  ( .D(N10338), .E(N10353), .CP(clk), .Q(
        \entry[4][21] ) );
  EDFQD1 \entry_reg[4][20]  ( .D(N10337), .E(N10353), .CP(clk), .Q(
        \entry[4][20] ) );
  EDFQD1 \entry_reg[4][19]  ( .D(N10336), .E(N10353), .CP(clk), .Q(
        \entry[4][19] ) );
  EDFQD1 \entry_reg[4][18]  ( .D(N10335), .E(N10353), .CP(clk), .Q(
        \entry[4][18] ) );
  EDFQD1 \entry_reg[4][17]  ( .D(N10334), .E(N10353), .CP(clk), .Q(
        \entry[4][17] ) );
  EDFQD1 \entry_reg[4][16]  ( .D(N10333), .E(N10353), .CP(clk), .Q(
        \entry[4][16] ) );
  EDFQD1 \entry_reg[4][15]  ( .D(N10332), .E(N10353), .CP(clk), .Q(
        \entry[4][15] ) );
  EDFQD1 \entry_reg[4][14]  ( .D(N10331), .E(N10353), .CP(clk), .Q(
        \entry[4][14] ) );
  EDFQD1 \entry_reg[4][13]  ( .D(N10330), .E(N10353), .CP(clk), .Q(
        \entry[4][13] ) );
  EDFQD1 \entry_reg[4][12]  ( .D(N10329), .E(N10353), .CP(clk), .Q(
        \entry[4][12] ) );
  EDFQD1 \entry_reg[4][11]  ( .D(N10328), .E(N10353), .CP(clk), .Q(
        \entry[4][11] ) );
  EDFQD1 \entry_reg[4][10]  ( .D(N10327), .E(N10353), .CP(clk), .Q(
        \entry[4][10] ) );
  EDFQD1 \entry_reg[4][9]  ( .D(N10326), .E(N10353), .CP(clk), .Q(
        \entry[4][9] ) );
  EDFQD1 \entry_reg[4][8]  ( .D(N10325), .E(N10353), .CP(clk), .Q(
        \entry[4][8] ) );
  EDFQD1 \entry_reg[4][7]  ( .D(N10324), .E(N10353), .CP(clk), .Q(
        \entry[4][7] ) );
  EDFQD1 \entry_reg[4][6]  ( .D(N10323), .E(N10353), .CP(clk), .Q(
        \entry[4][6] ) );
  EDFQD1 \entry_reg[4][5]  ( .D(N10322), .E(N10353), .CP(clk), .Q(
        \entry[4][5] ) );
  EDFQD1 \entry_reg[4][4]  ( .D(N10321), .E(N10353), .CP(clk), .Q(
        \entry[4][4] ) );
  EDFQD1 \entry_reg[4][3]  ( .D(N10320), .E(N10353), .CP(clk), .Q(
        \entry[4][3] ) );
  EDFQD1 \entry_reg[4][2]  ( .D(N10319), .E(N10353), .CP(clk), .Q(
        \entry[4][2] ) );
  EDFQD1 \entry_reg[4][1]  ( .D(N10318), .E(N10353), .CP(clk), .Q(
        \entry[4][1] ) );
  EDFQD1 \entry_reg[4][0]  ( .D(N10317), .E(N10353), .CP(clk), .Q(
        \entry[4][0] ) );
  EDFQD1 \entry_reg[3][31]  ( .D(N10348), .E(N10352), .CP(clk), .Q(
        \entry[3][31] ) );
  EDFQD1 \entry_reg[3][30]  ( .D(N10347), .E(N10352), .CP(clk), .Q(
        \entry[3][30] ) );
  EDFQD1 \entry_reg[3][29]  ( .D(N10346), .E(N10352), .CP(clk), .Q(
        \entry[3][29] ) );
  EDFQD1 \entry_reg[3][28]  ( .D(N10345), .E(N10352), .CP(clk), .Q(
        \entry[3][28] ) );
  EDFQD1 \entry_reg[3][27]  ( .D(N10344), .E(N10352), .CP(clk), .Q(
        \entry[3][27] ) );
  EDFQD1 \entry_reg[3][26]  ( .D(N10343), .E(N10352), .CP(clk), .Q(
        \entry[3][26] ) );
  EDFQD1 \entry_reg[3][25]  ( .D(N10342), .E(N10352), .CP(clk), .Q(
        \entry[3][25] ) );
  EDFQD1 \entry_reg[3][24]  ( .D(N10341), .E(N10352), .CP(clk), .Q(
        \entry[3][24] ) );
  EDFQD1 \entry_reg[3][23]  ( .D(N10340), .E(N10352), .CP(clk), .Q(
        \entry[3][23] ) );
  EDFQD1 \entry_reg[3][22]  ( .D(N10339), .E(N10352), .CP(clk), .Q(
        \entry[3][22] ) );
  EDFQD1 \entry_reg[3][21]  ( .D(N10338), .E(N10352), .CP(clk), .Q(
        \entry[3][21] ) );
  EDFQD1 \entry_reg[3][20]  ( .D(N10337), .E(N10352), .CP(clk), .Q(
        \entry[3][20] ) );
  EDFQD1 \entry_reg[3][19]  ( .D(N10336), .E(N10352), .CP(clk), .Q(
        \entry[3][19] ) );
  EDFQD1 \entry_reg[3][18]  ( .D(N10335), .E(N10352), .CP(clk), .Q(
        \entry[3][18] ) );
  EDFQD1 \entry_reg[3][17]  ( .D(N10334), .E(N10352), .CP(clk), .Q(
        \entry[3][17] ) );
  EDFQD1 \entry_reg[3][16]  ( .D(N10333), .E(N10352), .CP(clk), .Q(
        \entry[3][16] ) );
  EDFQD1 \entry_reg[3][15]  ( .D(N10332), .E(N10352), .CP(clk), .Q(
        \entry[3][15] ) );
  EDFQD1 \entry_reg[3][14]  ( .D(N10331), .E(N10352), .CP(clk), .Q(
        \entry[3][14] ) );
  EDFQD1 \entry_reg[3][13]  ( .D(N10330), .E(N10352), .CP(clk), .Q(
        \entry[3][13] ) );
  EDFQD1 \entry_reg[3][12]  ( .D(N10329), .E(N10352), .CP(clk), .Q(
        \entry[3][12] ) );
  EDFQD1 \entry_reg[3][11]  ( .D(N10328), .E(N10352), .CP(clk), .Q(
        \entry[3][11] ) );
  EDFQD1 \entry_reg[3][10]  ( .D(N10327), .E(N10352), .CP(clk), .Q(
        \entry[3][10] ) );
  EDFQD1 \entry_reg[3][9]  ( .D(N10326), .E(N10352), .CP(clk), .Q(
        \entry[3][9] ) );
  EDFQD1 \entry_reg[3][8]  ( .D(N10325), .E(N10352), .CP(clk), .Q(
        \entry[3][8] ) );
  EDFQD1 \entry_reg[3][7]  ( .D(N10324), .E(N10352), .CP(clk), .Q(
        \entry[3][7] ) );
  EDFQD1 \entry_reg[3][6]  ( .D(N10323), .E(N10352), .CP(clk), .Q(
        \entry[3][6] ) );
  EDFQD1 \entry_reg[3][5]  ( .D(N10322), .E(N10352), .CP(clk), .Q(
        \entry[3][5] ) );
  EDFQD1 \entry_reg[3][4]  ( .D(N10321), .E(N10352), .CP(clk), .Q(
        \entry[3][4] ) );
  EDFQD1 \entry_reg[3][3]  ( .D(N10320), .E(N10352), .CP(clk), .Q(
        \entry[3][3] ) );
  EDFQD1 \entry_reg[3][2]  ( .D(N10319), .E(N10352), .CP(clk), .Q(
        \entry[3][2] ) );
  EDFQD1 \entry_reg[3][1]  ( .D(N10318), .E(N10352), .CP(clk), .Q(
        \entry[3][1] ) );
  EDFQD1 \entry_reg[3][0]  ( .D(N10317), .E(N10352), .CP(clk), .Q(
        \entry[3][0] ) );
  EDFQD1 \entry_reg[2][31]  ( .D(N10348), .E(N10351), .CP(clk), .Q(
        \entry[2][31] ) );
  EDFQD1 \entry_reg[2][30]  ( .D(N10347), .E(N10351), .CP(clk), .Q(
        \entry[2][30] ) );
  EDFQD1 \entry_reg[2][29]  ( .D(N10346), .E(N10351), .CP(clk), .Q(
        \entry[2][29] ) );
  EDFQD1 \entry_reg[2][28]  ( .D(N10345), .E(N10351), .CP(clk), .Q(
        \entry[2][28] ) );
  EDFQD1 \entry_reg[2][27]  ( .D(N10344), .E(N10351), .CP(clk), .Q(
        \entry[2][27] ) );
  EDFQD1 \entry_reg[2][26]  ( .D(N10343), .E(N10351), .CP(clk), .Q(
        \entry[2][26] ) );
  EDFQD1 \entry_reg[2][25]  ( .D(N10342), .E(N10351), .CP(clk), .Q(
        \entry[2][25] ) );
  EDFQD1 \entry_reg[2][24]  ( .D(N10341), .E(N10351), .CP(clk), .Q(
        \entry[2][24] ) );
  EDFQD1 \entry_reg[2][23]  ( .D(N10340), .E(N10351), .CP(clk), .Q(
        \entry[2][23] ) );
  EDFQD1 \entry_reg[2][22]  ( .D(N10339), .E(N10351), .CP(clk), .Q(
        \entry[2][22] ) );
  EDFQD1 \entry_reg[2][21]  ( .D(N10338), .E(N10351), .CP(clk), .Q(
        \entry[2][21] ) );
  EDFQD1 \entry_reg[2][20]  ( .D(N10337), .E(N10351), .CP(clk), .Q(
        \entry[2][20] ) );
  EDFQD1 \entry_reg[2][19]  ( .D(N10336), .E(N10351), .CP(clk), .Q(
        \entry[2][19] ) );
  EDFQD1 \entry_reg[2][18]  ( .D(N10335), .E(N10351), .CP(clk), .Q(
        \entry[2][18] ) );
  EDFQD1 \entry_reg[2][17]  ( .D(N10334), .E(N10351), .CP(clk), .Q(
        \entry[2][17] ) );
  EDFQD1 \entry_reg[2][16]  ( .D(N10333), .E(N10351), .CP(clk), .Q(
        \entry[2][16] ) );
  EDFQD1 \entry_reg[2][15]  ( .D(N10332), .E(N10351), .CP(clk), .Q(
        \entry[2][15] ) );
  EDFQD1 \entry_reg[2][14]  ( .D(N10331), .E(N10351), .CP(clk), .Q(
        \entry[2][14] ) );
  EDFQD1 \entry_reg[2][13]  ( .D(N10330), .E(N10351), .CP(clk), .Q(
        \entry[2][13] ) );
  EDFQD1 \entry_reg[2][12]  ( .D(N10329), .E(N10351), .CP(clk), .Q(
        \entry[2][12] ) );
  EDFQD1 \entry_reg[2][11]  ( .D(N10328), .E(N10351), .CP(clk), .Q(
        \entry[2][11] ) );
  EDFQD1 \entry_reg[2][10]  ( .D(N10327), .E(N10351), .CP(clk), .Q(
        \entry[2][10] ) );
  EDFQD1 \entry_reg[2][9]  ( .D(N10326), .E(N10351), .CP(clk), .Q(
        \entry[2][9] ) );
  EDFQD1 \entry_reg[2][8]  ( .D(N10325), .E(N10351), .CP(clk), .Q(
        \entry[2][8] ) );
  EDFQD1 \entry_reg[2][7]  ( .D(N10324), .E(N10351), .CP(clk), .Q(
        \entry[2][7] ) );
  EDFQD1 \entry_reg[2][6]  ( .D(N10323), .E(N10351), .CP(clk), .Q(
        \entry[2][6] ) );
  EDFQD1 \entry_reg[2][5]  ( .D(N10322), .E(N10351), .CP(clk), .Q(
        \entry[2][5] ) );
  EDFQD1 \entry_reg[2][4]  ( .D(N10321), .E(N10351), .CP(clk), .Q(
        \entry[2][4] ) );
  EDFQD1 \entry_reg[2][3]  ( .D(N10320), .E(N10351), .CP(clk), .Q(
        \entry[2][3] ) );
  EDFQD1 \entry_reg[2][2]  ( .D(N10319), .E(N10351), .CP(clk), .Q(
        \entry[2][2] ) );
  EDFQD1 \entry_reg[2][1]  ( .D(N10318), .E(N10351), .CP(clk), .Q(
        \entry[2][1] ) );
  EDFQD1 \entry_reg[2][0]  ( .D(N10317), .E(N10351), .CP(clk), .Q(
        \entry[2][0] ) );
  EDFQD1 \entry_reg[1][31]  ( .D(N10348), .E(N10350), .CP(clk), .Q(
        \entry[1][31] ) );
  EDFQD1 \entry_reg[1][30]  ( .D(N10347), .E(N10350), .CP(clk), .Q(
        \entry[1][30] ) );
  EDFQD1 \entry_reg[1][29]  ( .D(N10346), .E(N10350), .CP(clk), .Q(
        \entry[1][29] ) );
  EDFQD1 \entry_reg[1][28]  ( .D(N10345), .E(N10350), .CP(clk), .Q(
        \entry[1][28] ) );
  EDFQD1 \entry_reg[1][27]  ( .D(N10344), .E(N10350), .CP(clk), .Q(
        \entry[1][27] ) );
  EDFQD1 \entry_reg[1][26]  ( .D(N10343), .E(N10350), .CP(clk), .Q(
        \entry[1][26] ) );
  EDFQD1 \entry_reg[1][25]  ( .D(N10342), .E(N10350), .CP(clk), .Q(
        \entry[1][25] ) );
  EDFQD1 \entry_reg[1][24]  ( .D(N10341), .E(N10350), .CP(clk), .Q(
        \entry[1][24] ) );
  EDFQD1 \entry_reg[1][23]  ( .D(N10340), .E(N10350), .CP(clk), .Q(
        \entry[1][23] ) );
  EDFQD1 \entry_reg[1][22]  ( .D(N10339), .E(N10350), .CP(clk), .Q(
        \entry[1][22] ) );
  EDFQD1 \entry_reg[1][21]  ( .D(N10338), .E(N10350), .CP(clk), .Q(
        \entry[1][21] ) );
  EDFQD1 \entry_reg[1][20]  ( .D(N10337), .E(N10350), .CP(clk), .Q(
        \entry[1][20] ) );
  EDFQD1 \entry_reg[1][19]  ( .D(N10336), .E(N10350), .CP(clk), .Q(
        \entry[1][19] ) );
  EDFQD1 \entry_reg[1][18]  ( .D(N10335), .E(N10350), .CP(clk), .Q(
        \entry[1][18] ) );
  EDFQD1 \entry_reg[1][17]  ( .D(N10334), .E(N10350), .CP(clk), .Q(
        \entry[1][17] ) );
  EDFQD1 \entry_reg[1][16]  ( .D(N10333), .E(N10350), .CP(clk), .Q(
        \entry[1][16] ) );
  EDFQD1 \entry_reg[1][15]  ( .D(N10332), .E(N10350), .CP(clk), .Q(
        \entry[1][15] ) );
  EDFQD1 \entry_reg[1][14]  ( .D(N10331), .E(N10350), .CP(clk), .Q(
        \entry[1][14] ) );
  EDFQD1 \entry_reg[1][13]  ( .D(N10330), .E(N10350), .CP(clk), .Q(
        \entry[1][13] ) );
  EDFQD1 \entry_reg[1][12]  ( .D(N10329), .E(N10350), .CP(clk), .Q(
        \entry[1][12] ) );
  EDFQD1 \entry_reg[1][11]  ( .D(N10328), .E(N10350), .CP(clk), .Q(
        \entry[1][11] ) );
  EDFQD1 \entry_reg[1][10]  ( .D(N10327), .E(N10350), .CP(clk), .Q(
        \entry[1][10] ) );
  EDFQD1 \entry_reg[1][9]  ( .D(N10326), .E(N10350), .CP(clk), .Q(
        \entry[1][9] ) );
  EDFQD1 \entry_reg[1][8]  ( .D(N10325), .E(N10350), .CP(clk), .Q(
        \entry[1][8] ) );
  EDFQD1 \entry_reg[1][7]  ( .D(N10324), .E(N10350), .CP(clk), .Q(
        \entry[1][7] ) );
  EDFQD1 \entry_reg[1][6]  ( .D(N10323), .E(N10350), .CP(clk), .Q(
        \entry[1][6] ) );
  EDFQD1 \entry_reg[1][5]  ( .D(N10322), .E(N10350), .CP(clk), .Q(
        \entry[1][5] ) );
  EDFQD1 \entry_reg[1][4]  ( .D(N10321), .E(N10350), .CP(clk), .Q(
        \entry[1][4] ) );
  EDFQD1 \entry_reg[1][3]  ( .D(N10320), .E(N10350), .CP(clk), .Q(
        \entry[1][3] ) );
  EDFQD1 \entry_reg[1][2]  ( .D(N10319), .E(N10350), .CP(clk), .Q(
        \entry[1][2] ) );
  EDFQD1 \entry_reg[1][1]  ( .D(N10318), .E(N10350), .CP(clk), .Q(
        \entry[1][1] ) );
  EDFQD1 \entry_reg[1][0]  ( .D(N10317), .E(N10350), .CP(clk), .Q(
        \entry[1][0] ) );
  EDFQD1 \entry_reg[0][31]  ( .D(N10348), .E(N10349), .CP(clk), .Q(
        \entry[0][31] ) );
  EDFQD1 \entry_reg[0][30]  ( .D(N10347), .E(N10349), .CP(clk), .Q(
        \entry[0][30] ) );
  EDFQD1 \entry_reg[0][29]  ( .D(N10346), .E(N10349), .CP(clk), .Q(
        \entry[0][29] ) );
  EDFQD1 \entry_reg[0][28]  ( .D(N10345), .E(N10349), .CP(clk), .Q(
        \entry[0][28] ) );
  EDFQD1 \entry_reg[0][27]  ( .D(N10344), .E(N10349), .CP(clk), .Q(
        \entry[0][27] ) );
  EDFQD1 \entry_reg[0][26]  ( .D(N10343), .E(N10349), .CP(clk), .Q(
        \entry[0][26] ) );
  EDFQD1 \entry_reg[0][25]  ( .D(N10342), .E(N10349), .CP(clk), .Q(
        \entry[0][25] ) );
  EDFQD1 \entry_reg[0][24]  ( .D(N10341), .E(N10349), .CP(clk), .Q(
        \entry[0][24] ) );
  EDFQD1 \entry_reg[0][23]  ( .D(N10340), .E(N10349), .CP(clk), .Q(
        \entry[0][23] ) );
  EDFQD1 \entry_reg[0][22]  ( .D(N10339), .E(N10349), .CP(clk), .Q(
        \entry[0][22] ) );
  EDFQD1 \entry_reg[0][21]  ( .D(N10338), .E(N10349), .CP(clk), .Q(
        \entry[0][21] ) );
  EDFQD1 \entry_reg[0][20]  ( .D(N10337), .E(N10349), .CP(clk), .Q(
        \entry[0][20] ) );
  EDFQD1 \entry_reg[0][19]  ( .D(N10336), .E(N10349), .CP(clk), .Q(
        \entry[0][19] ) );
  EDFQD1 \entry_reg[0][18]  ( .D(N10335), .E(N10349), .CP(clk), .Q(
        \entry[0][18] ) );
  EDFQD1 \entry_reg[0][17]  ( .D(N10334), .E(N10349), .CP(clk), .Q(
        \entry[0][17] ) );
  EDFQD1 \entry_reg[0][16]  ( .D(N10333), .E(N10349), .CP(clk), .Q(
        \entry[0][16] ) );
  EDFQD1 \entry_reg[0][15]  ( .D(N10332), .E(N10349), .CP(clk), .Q(
        \entry[0][15] ) );
  EDFQD1 \entry_reg[0][14]  ( .D(N10331), .E(N10349), .CP(clk), .Q(
        \entry[0][14] ) );
  EDFQD1 \entry_reg[0][13]  ( .D(N10330), .E(N10349), .CP(clk), .Q(
        \entry[0][13] ) );
  EDFQD1 \entry_reg[0][12]  ( .D(N10329), .E(N10349), .CP(clk), .Q(
        \entry[0][12] ) );
  EDFQD1 \entry_reg[0][11]  ( .D(N10328), .E(N10349), .CP(clk), .Q(
        \entry[0][11] ) );
  EDFQD1 \entry_reg[0][10]  ( .D(N10327), .E(N10349), .CP(clk), .Q(
        \entry[0][10] ) );
  EDFQD1 \entry_reg[0][9]  ( .D(N10326), .E(N10349), .CP(clk), .Q(
        \entry[0][9] ) );
  EDFQD1 \entry_reg[0][8]  ( .D(N10325), .E(N10349), .CP(clk), .Q(
        \entry[0][8] ) );
  EDFQD1 \entry_reg[0][7]  ( .D(N10324), .E(N10349), .CP(clk), .Q(
        \entry[0][7] ) );
  EDFQD1 \entry_reg[0][6]  ( .D(N10323), .E(N10349), .CP(clk), .Q(
        \entry[0][6] ) );
  EDFQD1 \entry_reg[0][5]  ( .D(N10322), .E(N10349), .CP(clk), .Q(
        \entry[0][5] ) );
  EDFQD1 \entry_reg[0][4]  ( .D(N10321), .E(N10349), .CP(clk), .Q(
        \entry[0][4] ) );
  EDFQD1 \entry_reg[0][3]  ( .D(N10320), .E(N10349), .CP(clk), .Q(
        \entry[0][3] ) );
  EDFQD1 \entry_reg[0][2]  ( .D(N10319), .E(N10349), .CP(clk), .Q(
        \entry[0][2] ) );
  EDFQD1 \entry_reg[0][1]  ( .D(N10318), .E(N10349), .CP(clk), .Q(
        \entry[0][1] ) );
  EDFQD1 \entry_reg[0][0]  ( .D(N10317), .E(N10349), .CP(clk), .Q(
        \entry[0][0] ) );
  OAI21D1 U2110 ( .A1(n3243), .A2(n3259), .B(n3260), .ZN(n3000) );
  OAI21D1 U2111 ( .A1(n3243), .A2(n3248), .B(n3249), .ZN(n2995) );
  OAI21D1 U2112 ( .A1(n3243), .A2(n3244), .B(n3245), .ZN(n2990) );
  OAI21D1 U2113 ( .A1(n3243), .A2(n3255), .B(n3256), .ZN(n2991) );
  OAI21D1 U2114 ( .A1(n3243), .A2(n3263), .B(n3264), .ZN(n2996) );
  OAI22D1 U2115 ( .A1(n3266), .A2(n3267), .B1(n3243), .B2(n3268), .ZN(n3005)
         );
  NR2D2 U2116 ( .A1(n2972), .A2(n2976), .ZN(N10352) );
  NR2D2 U2117 ( .A1(n2968), .A2(n2971), .ZN(N10362) );
  OAI21D1 U2118 ( .A1(n3243), .A2(n3250), .B(n3251), .ZN(n2994) );
  NR2D2 U2119 ( .A1(n2969), .A2(n2976), .ZN(N10356) );
  NR2D2 U2120 ( .A1(n2968), .A2(n2973), .ZN(N10358) );
  NR2D2 U2121 ( .A1(n2970), .A2(n2972), .ZN(N10359) );
  OAI21D1 U2122 ( .A1(n3243), .A2(n3261), .B(n3262), .ZN(n2999) );
  NR2D2 U2123 ( .A1(n2973), .A2(n2976), .ZN(N10350) );
  NR2D2 U2124 ( .A1(n2968), .A2(n2969), .ZN(N10364) );
  NR2D2 U2125 ( .A1(n2970), .A2(n2971), .ZN(N10361) );
  OAI22D1 U2126 ( .A1(n3244), .A2(n3270), .B1(n3316), .B2(n3338), .ZN(n3004)
         );
  OAI21D1 U2127 ( .A1(n3243), .A2(n3252), .B(n3253), .ZN(n2992) );
  NR2D2 U2128 ( .A1(n2969), .A2(n2977), .ZN(N10355) );
  NR2D2 U2129 ( .A1(n2971), .A2(n2976), .ZN(N10354) );
  NR2D2 U2130 ( .A1(n2968), .A2(n2972), .ZN(N10360) );
  NR2D2 U2131 ( .A1(n2970), .A2(n2973), .ZN(N10357) );
  OAI22D1 U2132 ( .A1(n3243), .A2(n3269), .B1(n3270), .B2(n3271), .ZN(n3002)
         );
  ND3D1 U2133 ( .A1(n3266), .A2(n3289), .A3(n3290), .ZN(n3271) );
  INR3D1 U2134 ( .A1(en), .B1(wr), .B2(rst), .ZN(N10366) );
  NR2D2 U2135 ( .A1(n2971), .A2(n2977), .ZN(N10353) );
  NR2D2 U2136 ( .A1(n2972), .A2(n2977), .ZN(N10351) );
  ND3D0 U2137 ( .A1(n2975), .A2(n2980), .A3(n2974), .ZN(n2977) );
  NR2D2 U2138 ( .A1(n2973), .A2(n2977), .ZN(N10349) );
  NR2D2 U2139 ( .A1(n2969), .A2(n2970), .ZN(N10363) );
  ND3D1 U2140 ( .A1(n2974), .A2(n2975), .A3(index[3]), .ZN(n2970) );
  TIEL U2141 ( .ZN(n2463) );
  ND3D0 U2142 ( .A1(index[0]), .A2(n2974), .A3(index[3]), .ZN(n2968) );
  CKND2D0 U2143 ( .A1(index[2]), .A2(index[1]), .ZN(n2969) );
  CKND2D0 U2144 ( .A1(index[2]), .A2(n2978), .ZN(n2971) );
  CKND2D0 U2145 ( .A1(index[1]), .A2(n2979), .ZN(n2972) );
  ND3D0 U2146 ( .A1(n2974), .A2(n2980), .A3(index[0]), .ZN(n2976) );
  AN3D0 U2147 ( .A1(n2981), .A2(en), .A3(wr), .Z(n2974) );
  CKND0 U2148 ( .I(index[3]), .ZN(n2980) );
  CKND0 U2149 ( .I(index[0]), .ZN(n2975) );
  CKND2D0 U2150 ( .A1(n2978), .A2(n2979), .ZN(n2973) );
  CKND0 U2151 ( .I(index[2]), .ZN(n2979) );
  CKND0 U2152 ( .I(index[1]), .ZN(n2978) );
  AN2D0 U2153 ( .A1(store_val[31]), .A2(n2981), .Z(N10348) );
  AN2D0 U2154 ( .A1(store_val[30]), .A2(n2981), .Z(N10347) );
  AN2D0 U2155 ( .A1(store_val[29]), .A2(n2981), .Z(N10346) );
  AN2D0 U2156 ( .A1(store_val[28]), .A2(n2981), .Z(N10345) );
  AN2D0 U2157 ( .A1(store_val[27]), .A2(n2981), .Z(N10344) );
  AN2D0 U2158 ( .A1(store_val[26]), .A2(n2981), .Z(N10343) );
  AN2D0 U2159 ( .A1(store_val[25]), .A2(n2981), .Z(N10342) );
  AN2D0 U2160 ( .A1(store_val[24]), .A2(n2981), .Z(N10341) );
  AN2D0 U2161 ( .A1(store_val[23]), .A2(n2981), .Z(N10340) );
  AN2D0 U2162 ( .A1(store_val[22]), .A2(n2981), .Z(N10339) );
  AN2D0 U2163 ( .A1(store_val[21]), .A2(n2981), .Z(N10338) );
  AN2D0 U2164 ( .A1(store_val[20]), .A2(n2981), .Z(N10337) );
  AN2D0 U2165 ( .A1(store_val[19]), .A2(n2981), .Z(N10336) );
  AN2D0 U2166 ( .A1(store_val[18]), .A2(n2981), .Z(N10335) );
  AN2D0 U2167 ( .A1(store_val[17]), .A2(n2981), .Z(N10334) );
  AN2D0 U2168 ( .A1(store_val[16]), .A2(n2981), .Z(N10333) );
  AN2D0 U2169 ( .A1(store_val[15]), .A2(n2981), .Z(N10332) );
  AN2D0 U2170 ( .A1(store_val[14]), .A2(n2981), .Z(N10331) );
  AN2D0 U2171 ( .A1(store_val[13]), .A2(n2981), .Z(N10330) );
  AN2D0 U2172 ( .A1(store_val[12]), .A2(n2981), .Z(N10329) );
  AN2D0 U2173 ( .A1(store_val[11]), .A2(n2981), .Z(N10328) );
  AN2D0 U2174 ( .A1(store_val[10]), .A2(n2981), .Z(N10327) );
  AN2D0 U2175 ( .A1(store_val[9]), .A2(n2981), .Z(N10326) );
  AN2D0 U2176 ( .A1(store_val[8]), .A2(n2981), .Z(N10325) );
  AN2D0 U2177 ( .A1(store_val[7]), .A2(n2981), .Z(N10324) );
  AN2D0 U2178 ( .A1(store_val[6]), .A2(n2981), .Z(N10323) );
  AN2D0 U2179 ( .A1(store_val[5]), .A2(n2981), .Z(N10322) );
  AN2D0 U2180 ( .A1(store_val[4]), .A2(n2981), .Z(N10321) );
  AN2D0 U2181 ( .A1(store_val[3]), .A2(n2981), .Z(N10320) );
  AN2D0 U2182 ( .A1(store_val[2]), .A2(n2981), .Z(N10319) );
  AN2D0 U2183 ( .A1(store_val[1]), .A2(n2981), .Z(N10318) );
  AN2D0 U2184 ( .A1(store_val[0]), .A2(n2981), .Z(N10317) );
  CKND0 U2185 ( .I(rst), .ZN(n2981) );
  ND4D0 U2186 ( .A1(n2982), .A2(n2983), .A3(n2984), .A4(n2985), .ZN(N10316) );
  AOI221D0 U2187 ( .A1(\entry[12][15] ), .A2(n2986), .B1(\entry[13][15] ), 
        .B2(n2987), .C(n2988), .ZN(n2985) );
  AO22D0 U2188 ( .A1(\entry[11][15] ), .A2(n2989), .B1(\entry[0][15] ), .B2(
        n2990), .Z(n2988) );
  AOI221D0 U2189 ( .A1(\entry[1][15] ), .A2(n2991), .B1(\entry[2][15] ), .B2(
        n2992), .C(n2993), .ZN(n2984) );
  AO22D0 U2190 ( .A1(\entry[4][15] ), .A2(n2994), .B1(\entry[3][15] ), .B2(
        n2995), .Z(n2993) );
  AOI221D0 U2191 ( .A1(\entry[7][15] ), .A2(n2996), .B1(\entry[10][15] ), .B2(
        n2997), .C(n2998), .ZN(n2983) );
  AO22D0 U2192 ( .A1(\entry[6][15] ), .A2(n2999), .B1(\entry[5][15] ), .B2(
        n3000), .Z(n2998) );
  AOI221D0 U2193 ( .A1(\entry[14][15] ), .A2(n3001), .B1(\entry[9][15] ), .B2(
        n3002), .C(n3003), .ZN(n2982) );
  AO22D0 U2194 ( .A1(\entry[15][15] ), .A2(n3004), .B1(\entry[8][15] ), .B2(
        n3005), .Z(n3003) );
  ND4D0 U2195 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .ZN(N10315) );
  AOI221D0 U2196 ( .A1(\entry[12][14] ), .A2(n2986), .B1(\entry[13][14] ), 
        .B2(n2987), .C(n3010), .ZN(n3009) );
  AO22D0 U2197 ( .A1(\entry[11][14] ), .A2(n2989), .B1(\entry[0][14] ), .B2(
        n2990), .Z(n3010) );
  AOI221D0 U2198 ( .A1(\entry[1][14] ), .A2(n2991), .B1(\entry[2][14] ), .B2(
        n2992), .C(n3011), .ZN(n3008) );
  AO22D0 U2199 ( .A1(\entry[4][14] ), .A2(n2994), .B1(\entry[3][14] ), .B2(
        n2995), .Z(n3011) );
  AOI221D0 U2200 ( .A1(\entry[7][14] ), .A2(n2996), .B1(\entry[10][14] ), .B2(
        n2997), .C(n3012), .ZN(n3007) );
  AO22D0 U2201 ( .A1(\entry[6][14] ), .A2(n2999), .B1(\entry[5][14] ), .B2(
        n3000), .Z(n3012) );
  AOI221D0 U2202 ( .A1(\entry[14][14] ), .A2(n3001), .B1(\entry[9][14] ), .B2(
        n3002), .C(n3013), .ZN(n3006) );
  AO22D0 U2203 ( .A1(\entry[15][14] ), .A2(n3004), .B1(\entry[8][14] ), .B2(
        n3005), .Z(n3013) );
  ND4D0 U2204 ( .A1(n3014), .A2(n3015), .A3(n3016), .A4(n3017), .ZN(N10314) );
  AOI221D0 U2205 ( .A1(\entry[12][13] ), .A2(n2986), .B1(\entry[13][13] ), 
        .B2(n2987), .C(n3018), .ZN(n3017) );
  AO22D0 U2206 ( .A1(\entry[11][13] ), .A2(n2989), .B1(\entry[0][13] ), .B2(
        n2990), .Z(n3018) );
  AOI221D0 U2207 ( .A1(\entry[1][13] ), .A2(n2991), .B1(\entry[2][13] ), .B2(
        n2992), .C(n3019), .ZN(n3016) );
  AO22D0 U2208 ( .A1(\entry[4][13] ), .A2(n2994), .B1(\entry[3][13] ), .B2(
        n2995), .Z(n3019) );
  AOI221D0 U2209 ( .A1(\entry[7][13] ), .A2(n2996), .B1(\entry[10][13] ), .B2(
        n2997), .C(n3020), .ZN(n3015) );
  AO22D0 U2210 ( .A1(\entry[6][13] ), .A2(n2999), .B1(\entry[5][13] ), .B2(
        n3000), .Z(n3020) );
  AOI221D0 U2211 ( .A1(\entry[14][13] ), .A2(n3001), .B1(\entry[9][13] ), .B2(
        n3002), .C(n3021), .ZN(n3014) );
  AO22D0 U2212 ( .A1(\entry[15][13] ), .A2(n3004), .B1(\entry[8][13] ), .B2(
        n3005), .Z(n3021) );
  ND4D0 U2213 ( .A1(n3022), .A2(n3023), .A3(n3024), .A4(n3025), .ZN(N10313) );
  AOI221D0 U2214 ( .A1(\entry[12][12] ), .A2(n2986), .B1(\entry[13][12] ), 
        .B2(n2987), .C(n3026), .ZN(n3025) );
  AO22D0 U2215 ( .A1(\entry[11][12] ), .A2(n2989), .B1(\entry[0][12] ), .B2(
        n2990), .Z(n3026) );
  AOI221D0 U2216 ( .A1(\entry[1][12] ), .A2(n2991), .B1(\entry[2][12] ), .B2(
        n2992), .C(n3027), .ZN(n3024) );
  AO22D0 U2217 ( .A1(\entry[4][12] ), .A2(n2994), .B1(\entry[3][12] ), .B2(
        n2995), .Z(n3027) );
  AOI221D0 U2218 ( .A1(\entry[7][12] ), .A2(n2996), .B1(\entry[10][12] ), .B2(
        n2997), .C(n3028), .ZN(n3023) );
  AO22D0 U2219 ( .A1(\entry[6][12] ), .A2(n2999), .B1(\entry[5][12] ), .B2(
        n3000), .Z(n3028) );
  AOI221D0 U2220 ( .A1(\entry[14][12] ), .A2(n3001), .B1(\entry[9][12] ), .B2(
        n3002), .C(n3029), .ZN(n3022) );
  AO22D0 U2221 ( .A1(\entry[15][12] ), .A2(n3004), .B1(\entry[8][12] ), .B2(
        n3005), .Z(n3029) );
  ND4D0 U2222 ( .A1(n3030), .A2(n3031), .A3(n3032), .A4(n3033), .ZN(N10312) );
  AOI221D0 U2223 ( .A1(\entry[12][11] ), .A2(n2986), .B1(\entry[13][11] ), 
        .B2(n2987), .C(n3034), .ZN(n3033) );
  AO22D0 U2224 ( .A1(\entry[11][11] ), .A2(n2989), .B1(\entry[0][11] ), .B2(
        n2990), .Z(n3034) );
  AOI221D0 U2225 ( .A1(\entry[1][11] ), .A2(n2991), .B1(\entry[2][11] ), .B2(
        n2992), .C(n3035), .ZN(n3032) );
  AO22D0 U2226 ( .A1(\entry[4][11] ), .A2(n2994), .B1(\entry[3][11] ), .B2(
        n2995), .Z(n3035) );
  AOI221D0 U2227 ( .A1(\entry[7][11] ), .A2(n2996), .B1(\entry[10][11] ), .B2(
        n2997), .C(n3036), .ZN(n3031) );
  AO22D0 U2228 ( .A1(\entry[6][11] ), .A2(n2999), .B1(\entry[5][11] ), .B2(
        n3000), .Z(n3036) );
  AOI221D0 U2229 ( .A1(\entry[14][11] ), .A2(n3001), .B1(\entry[9][11] ), .B2(
        n3002), .C(n3037), .ZN(n3030) );
  AO22D0 U2230 ( .A1(\entry[15][11] ), .A2(n3004), .B1(\entry[8][11] ), .B2(
        n3005), .Z(n3037) );
  ND4D0 U2231 ( .A1(n3038), .A2(n3039), .A3(n3040), .A4(n3041), .ZN(N10311) );
  AOI221D0 U2232 ( .A1(\entry[12][10] ), .A2(n2986), .B1(\entry[13][10] ), 
        .B2(n2987), .C(n3042), .ZN(n3041) );
  AO22D0 U2233 ( .A1(\entry[11][10] ), .A2(n2989), .B1(\entry[0][10] ), .B2(
        n2990), .Z(n3042) );
  AOI221D0 U2234 ( .A1(\entry[1][10] ), .A2(n2991), .B1(\entry[2][10] ), .B2(
        n2992), .C(n3043), .ZN(n3040) );
  AO22D0 U2235 ( .A1(\entry[4][10] ), .A2(n2994), .B1(\entry[3][10] ), .B2(
        n2995), .Z(n3043) );
  AOI221D0 U2236 ( .A1(\entry[7][10] ), .A2(n2996), .B1(\entry[10][10] ), .B2(
        n2997), .C(n3044), .ZN(n3039) );
  AO22D0 U2237 ( .A1(\entry[6][10] ), .A2(n2999), .B1(\entry[5][10] ), .B2(
        n3000), .Z(n3044) );
  AOI221D0 U2238 ( .A1(\entry[14][10] ), .A2(n3001), .B1(\entry[9][10] ), .B2(
        n3002), .C(n3045), .ZN(n3038) );
  AO22D0 U2239 ( .A1(\entry[15][10] ), .A2(n3004), .B1(\entry[8][10] ), .B2(
        n3005), .Z(n3045) );
  ND4D0 U2240 ( .A1(n3046), .A2(n3047), .A3(n3048), .A4(n3049), .ZN(N10310) );
  AOI221D0 U2241 ( .A1(\entry[12][9] ), .A2(n2986), .B1(\entry[13][9] ), .B2(
        n2987), .C(n3050), .ZN(n3049) );
  AO22D0 U2242 ( .A1(\entry[11][9] ), .A2(n2989), .B1(\entry[0][9] ), .B2(
        n2990), .Z(n3050) );
  AOI221D0 U2243 ( .A1(\entry[1][9] ), .A2(n2991), .B1(\entry[2][9] ), .B2(
        n2992), .C(n3051), .ZN(n3048) );
  AO22D0 U2244 ( .A1(\entry[4][9] ), .A2(n2994), .B1(\entry[3][9] ), .B2(n2995), .Z(n3051) );
  AOI221D0 U2245 ( .A1(\entry[7][9] ), .A2(n2996), .B1(\entry[10][9] ), .B2(
        n2997), .C(n3052), .ZN(n3047) );
  AO22D0 U2246 ( .A1(\entry[6][9] ), .A2(n2999), .B1(\entry[5][9] ), .B2(n3000), .Z(n3052) );
  AOI221D0 U2247 ( .A1(\entry[14][9] ), .A2(n3001), .B1(\entry[9][9] ), .B2(
        n3002), .C(n3053), .ZN(n3046) );
  AO22D0 U2248 ( .A1(\entry[15][9] ), .A2(n3004), .B1(\entry[8][9] ), .B2(
        n3005), .Z(n3053) );
  ND4D0 U2249 ( .A1(n3054), .A2(n3055), .A3(n3056), .A4(n3057), .ZN(N10309) );
  AOI221D0 U2250 ( .A1(\entry[12][8] ), .A2(n2986), .B1(\entry[13][8] ), .B2(
        n2987), .C(n3058), .ZN(n3057) );
  AO22D0 U2251 ( .A1(\entry[11][8] ), .A2(n2989), .B1(\entry[0][8] ), .B2(
        n2990), .Z(n3058) );
  AOI221D0 U2252 ( .A1(\entry[1][8] ), .A2(n2991), .B1(\entry[2][8] ), .B2(
        n2992), .C(n3059), .ZN(n3056) );
  AO22D0 U2253 ( .A1(\entry[4][8] ), .A2(n2994), .B1(\entry[3][8] ), .B2(n2995), .Z(n3059) );
  AOI221D0 U2254 ( .A1(\entry[7][8] ), .A2(n2996), .B1(\entry[10][8] ), .B2(
        n2997), .C(n3060), .ZN(n3055) );
  AO22D0 U2255 ( .A1(\entry[6][8] ), .A2(n2999), .B1(\entry[5][8] ), .B2(n3000), .Z(n3060) );
  AOI221D0 U2256 ( .A1(\entry[14][8] ), .A2(n3001), .B1(\entry[9][8] ), .B2(
        n3002), .C(n3061), .ZN(n3054) );
  AO22D0 U2257 ( .A1(\entry[15][8] ), .A2(n3004), .B1(\entry[8][8] ), .B2(
        n3005), .Z(n3061) );
  ND4D0 U2258 ( .A1(n3062), .A2(n3063), .A3(n3064), .A4(n3065), .ZN(N10308) );
  AOI221D0 U2259 ( .A1(\entry[12][7] ), .A2(n2986), .B1(\entry[13][7] ), .B2(
        n2987), .C(n3066), .ZN(n3065) );
  AO22D0 U2260 ( .A1(\entry[11][7] ), .A2(n2989), .B1(\entry[0][7] ), .B2(
        n2990), .Z(n3066) );
  AOI221D0 U2261 ( .A1(\entry[1][7] ), .A2(n2991), .B1(\entry[2][7] ), .B2(
        n2992), .C(n3067), .ZN(n3064) );
  AO22D0 U2262 ( .A1(\entry[4][7] ), .A2(n2994), .B1(\entry[3][7] ), .B2(n2995), .Z(n3067) );
  AOI221D0 U2263 ( .A1(\entry[7][7] ), .A2(n2996), .B1(\entry[10][7] ), .B2(
        n2997), .C(n3068), .ZN(n3063) );
  AO22D0 U2264 ( .A1(\entry[6][7] ), .A2(n2999), .B1(\entry[5][7] ), .B2(n3000), .Z(n3068) );
  AOI221D0 U2265 ( .A1(\entry[14][7] ), .A2(n3001), .B1(\entry[9][7] ), .B2(
        n3002), .C(n3069), .ZN(n3062) );
  AO22D0 U2266 ( .A1(\entry[15][7] ), .A2(n3004), .B1(\entry[8][7] ), .B2(
        n3005), .Z(n3069) );
  ND4D0 U2267 ( .A1(n3070), .A2(n3071), .A3(n3072), .A4(n3073), .ZN(N10307) );
  AOI221D0 U2268 ( .A1(\entry[12][6] ), .A2(n2986), .B1(\entry[13][6] ), .B2(
        n2987), .C(n3074), .ZN(n3073) );
  AO22D0 U2269 ( .A1(\entry[11][6] ), .A2(n2989), .B1(\entry[0][6] ), .B2(
        n2990), .Z(n3074) );
  AOI221D0 U2270 ( .A1(\entry[1][6] ), .A2(n2991), .B1(\entry[2][6] ), .B2(
        n2992), .C(n3075), .ZN(n3072) );
  AO22D0 U2271 ( .A1(\entry[4][6] ), .A2(n2994), .B1(\entry[3][6] ), .B2(n2995), .Z(n3075) );
  AOI221D0 U2272 ( .A1(\entry[7][6] ), .A2(n2996), .B1(\entry[10][6] ), .B2(
        n2997), .C(n3076), .ZN(n3071) );
  AO22D0 U2273 ( .A1(\entry[6][6] ), .A2(n2999), .B1(\entry[5][6] ), .B2(n3000), .Z(n3076) );
  AOI221D0 U2274 ( .A1(\entry[14][6] ), .A2(n3001), .B1(\entry[9][6] ), .B2(
        n3002), .C(n3077), .ZN(n3070) );
  AO22D0 U2275 ( .A1(\entry[15][6] ), .A2(n3004), .B1(\entry[8][6] ), .B2(
        n3005), .Z(n3077) );
  ND4D0 U2276 ( .A1(n3078), .A2(n3079), .A3(n3080), .A4(n3081), .ZN(N10306) );
  AOI221D0 U2277 ( .A1(\entry[12][5] ), .A2(n2986), .B1(\entry[13][5] ), .B2(
        n2987), .C(n3082), .ZN(n3081) );
  AO22D0 U2278 ( .A1(\entry[11][5] ), .A2(n2989), .B1(\entry[0][5] ), .B2(
        n2990), .Z(n3082) );
  AOI221D0 U2279 ( .A1(\entry[1][5] ), .A2(n2991), .B1(\entry[2][5] ), .B2(
        n2992), .C(n3083), .ZN(n3080) );
  AO22D0 U2280 ( .A1(\entry[4][5] ), .A2(n2994), .B1(\entry[3][5] ), .B2(n2995), .Z(n3083) );
  AOI221D0 U2281 ( .A1(\entry[7][5] ), .A2(n2996), .B1(\entry[10][5] ), .B2(
        n2997), .C(n3084), .ZN(n3079) );
  AO22D0 U2282 ( .A1(\entry[6][5] ), .A2(n2999), .B1(\entry[5][5] ), .B2(n3000), .Z(n3084) );
  AOI221D0 U2283 ( .A1(\entry[14][5] ), .A2(n3001), .B1(\entry[9][5] ), .B2(
        n3002), .C(n3085), .ZN(n3078) );
  AO22D0 U2284 ( .A1(\entry[15][5] ), .A2(n3004), .B1(\entry[8][5] ), .B2(
        n3005), .Z(n3085) );
  ND4D0 U2285 ( .A1(n3086), .A2(n3087), .A3(n3088), .A4(n3089), .ZN(N10305) );
  AOI221D0 U2286 ( .A1(\entry[12][4] ), .A2(n2986), .B1(\entry[13][4] ), .B2(
        n2987), .C(n3090), .ZN(n3089) );
  AO22D0 U2287 ( .A1(\entry[11][4] ), .A2(n2989), .B1(\entry[0][4] ), .B2(
        n2990), .Z(n3090) );
  AOI221D0 U2288 ( .A1(\entry[1][4] ), .A2(n2991), .B1(\entry[2][4] ), .B2(
        n2992), .C(n3091), .ZN(n3088) );
  AO22D0 U2289 ( .A1(\entry[4][4] ), .A2(n2994), .B1(\entry[3][4] ), .B2(n2995), .Z(n3091) );
  AOI221D0 U2290 ( .A1(\entry[7][4] ), .A2(n2996), .B1(\entry[10][4] ), .B2(
        n2997), .C(n3092), .ZN(n3087) );
  AO22D0 U2291 ( .A1(\entry[6][4] ), .A2(n2999), .B1(\entry[5][4] ), .B2(n3000), .Z(n3092) );
  AOI221D0 U2292 ( .A1(\entry[14][4] ), .A2(n3001), .B1(\entry[9][4] ), .B2(
        n3002), .C(n3093), .ZN(n3086) );
  AO22D0 U2293 ( .A1(\entry[15][4] ), .A2(n3004), .B1(\entry[8][4] ), .B2(
        n3005), .Z(n3093) );
  ND4D0 U2294 ( .A1(n3094), .A2(n3095), .A3(n3096), .A4(n3097), .ZN(N10304) );
  AOI221D0 U2295 ( .A1(\entry[12][3] ), .A2(n2986), .B1(\entry[13][3] ), .B2(
        n2987), .C(n3098), .ZN(n3097) );
  AO22D0 U2296 ( .A1(\entry[11][3] ), .A2(n2989), .B1(\entry[0][3] ), .B2(
        n2990), .Z(n3098) );
  AOI221D0 U2297 ( .A1(\entry[1][3] ), .A2(n2991), .B1(\entry[2][3] ), .B2(
        n2992), .C(n3099), .ZN(n3096) );
  AO22D0 U2298 ( .A1(\entry[4][3] ), .A2(n2994), .B1(\entry[3][3] ), .B2(n2995), .Z(n3099) );
  AOI221D0 U2299 ( .A1(\entry[7][3] ), .A2(n2996), .B1(\entry[10][3] ), .B2(
        n2997), .C(n3100), .ZN(n3095) );
  AO22D0 U2300 ( .A1(\entry[6][3] ), .A2(n2999), .B1(\entry[5][3] ), .B2(n3000), .Z(n3100) );
  AOI221D0 U2301 ( .A1(\entry[14][3] ), .A2(n3001), .B1(\entry[9][3] ), .B2(
        n3002), .C(n3101), .ZN(n3094) );
  AO22D0 U2302 ( .A1(\entry[15][3] ), .A2(n3004), .B1(\entry[8][3] ), .B2(
        n3005), .Z(n3101) );
  ND4D0 U2303 ( .A1(n3102), .A2(n3103), .A3(n3104), .A4(n3105), .ZN(N10303) );
  AOI221D0 U2304 ( .A1(\entry[12][2] ), .A2(n2986), .B1(\entry[13][2] ), .B2(
        n2987), .C(n3106), .ZN(n3105) );
  AO22D0 U2305 ( .A1(\entry[11][2] ), .A2(n2989), .B1(\entry[0][2] ), .B2(
        n2990), .Z(n3106) );
  AOI221D0 U2306 ( .A1(\entry[1][2] ), .A2(n2991), .B1(\entry[2][2] ), .B2(
        n2992), .C(n3107), .ZN(n3104) );
  AO22D0 U2307 ( .A1(\entry[4][2] ), .A2(n2994), .B1(\entry[3][2] ), .B2(n2995), .Z(n3107) );
  AOI221D0 U2308 ( .A1(\entry[7][2] ), .A2(n2996), .B1(\entry[10][2] ), .B2(
        n2997), .C(n3108), .ZN(n3103) );
  AO22D0 U2309 ( .A1(\entry[6][2] ), .A2(n2999), .B1(\entry[5][2] ), .B2(n3000), .Z(n3108) );
  AOI221D0 U2310 ( .A1(\entry[14][2] ), .A2(n3001), .B1(\entry[9][2] ), .B2(
        n3002), .C(n3109), .ZN(n3102) );
  AO22D0 U2311 ( .A1(\entry[15][2] ), .A2(n3004), .B1(\entry[8][2] ), .B2(
        n3005), .Z(n3109) );
  ND4D0 U2312 ( .A1(n3110), .A2(n3111), .A3(n3112), .A4(n3113), .ZN(N10302) );
  AOI221D0 U2313 ( .A1(\entry[12][1] ), .A2(n2986), .B1(\entry[13][1] ), .B2(
        n2987), .C(n3114), .ZN(n3113) );
  AO22D0 U2314 ( .A1(\entry[11][1] ), .A2(n2989), .B1(\entry[0][1] ), .B2(
        n2990), .Z(n3114) );
  AOI221D0 U2315 ( .A1(\entry[1][1] ), .A2(n2991), .B1(\entry[2][1] ), .B2(
        n2992), .C(n3115), .ZN(n3112) );
  AO22D0 U2316 ( .A1(\entry[4][1] ), .A2(n2994), .B1(\entry[3][1] ), .B2(n2995), .Z(n3115) );
  AOI221D0 U2317 ( .A1(\entry[7][1] ), .A2(n2996), .B1(\entry[10][1] ), .B2(
        n2997), .C(n3116), .ZN(n3111) );
  AO22D0 U2318 ( .A1(\entry[6][1] ), .A2(n2999), .B1(\entry[5][1] ), .B2(n3000), .Z(n3116) );
  AOI221D0 U2319 ( .A1(\entry[14][1] ), .A2(n3001), .B1(\entry[9][1] ), .B2(
        n3002), .C(n3117), .ZN(n3110) );
  AO22D0 U2320 ( .A1(\entry[15][1] ), .A2(n3004), .B1(\entry[8][1] ), .B2(
        n3005), .Z(n3117) );
  ND4D0 U2321 ( .A1(n3118), .A2(n3119), .A3(n3120), .A4(n3121), .ZN(N10301) );
  AOI221D0 U2322 ( .A1(\entry[12][0] ), .A2(n2986), .B1(\entry[13][0] ), .B2(
        n2987), .C(n3122), .ZN(n3121) );
  AO22D0 U2323 ( .A1(\entry[11][0] ), .A2(n2989), .B1(\entry[0][0] ), .B2(
        n2990), .Z(n3122) );
  AOI221D0 U2324 ( .A1(\entry[1][0] ), .A2(n2991), .B1(\entry[2][0] ), .B2(
        n2992), .C(n3123), .ZN(n3120) );
  AO22D0 U2325 ( .A1(\entry[4][0] ), .A2(n2994), .B1(\entry[3][0] ), .B2(n2995), .Z(n3123) );
  AOI221D0 U2326 ( .A1(\entry[7][0] ), .A2(n2996), .B1(\entry[10][0] ), .B2(
        n2997), .C(n3124), .ZN(n3119) );
  AO22D0 U2327 ( .A1(\entry[6][0] ), .A2(n2999), .B1(\entry[5][0] ), .B2(n3000), .Z(n3124) );
  AOI221D0 U2328 ( .A1(\entry[14][0] ), .A2(n3001), .B1(\entry[9][0] ), .B2(
        n3002), .C(n3125), .ZN(n3118) );
  AO22D0 U2329 ( .A1(\entry[15][0] ), .A2(n3004), .B1(\entry[8][0] ), .B2(
        n3005), .Z(n3125) );
  ND4D0 U2330 ( .A1(n3126), .A2(n3127), .A3(n3128), .A4(n3129), .ZN(N10299) );
  AOI221D0 U2331 ( .A1(\entry[12][31] ), .A2(n2986), .B1(\entry[13][31] ), 
        .B2(n2987), .C(n3130), .ZN(n3129) );
  AO22D0 U2332 ( .A1(\entry[11][31] ), .A2(n2989), .B1(\entry[0][31] ), .B2(
        n2990), .Z(n3130) );
  AOI221D0 U2333 ( .A1(\entry[1][31] ), .A2(n2991), .B1(\entry[2][31] ), .B2(
        n2992), .C(n3131), .ZN(n3128) );
  AO22D0 U2334 ( .A1(\entry[4][31] ), .A2(n2994), .B1(\entry[3][31] ), .B2(
        n2995), .Z(n3131) );
  AOI221D0 U2335 ( .A1(\entry[7][31] ), .A2(n2996), .B1(\entry[10][31] ), .B2(
        n2997), .C(n3132), .ZN(n3127) );
  AO22D0 U2336 ( .A1(\entry[6][31] ), .A2(n2999), .B1(\entry[5][31] ), .B2(
        n3000), .Z(n3132) );
  AOI221D0 U2337 ( .A1(\entry[14][31] ), .A2(n3001), .B1(\entry[9][31] ), .B2(
        n3002), .C(n3133), .ZN(n3126) );
  AO22D0 U2338 ( .A1(\entry[15][31] ), .A2(n3004), .B1(\entry[8][31] ), .B2(
        n3005), .Z(n3133) );
  ND4D0 U2339 ( .A1(n3134), .A2(n3135), .A3(n3136), .A4(n3137), .ZN(N10298) );
  AOI221D0 U2340 ( .A1(\entry[12][30] ), .A2(n2986), .B1(\entry[13][30] ), 
        .B2(n2987), .C(n3138), .ZN(n3137) );
  AO22D0 U2341 ( .A1(\entry[11][30] ), .A2(n2989), .B1(\entry[0][30] ), .B2(
        n2990), .Z(n3138) );
  AOI221D0 U2342 ( .A1(\entry[1][30] ), .A2(n2991), .B1(\entry[2][30] ), .B2(
        n2992), .C(n3139), .ZN(n3136) );
  AO22D0 U2343 ( .A1(\entry[4][30] ), .A2(n2994), .B1(\entry[3][30] ), .B2(
        n2995), .Z(n3139) );
  AOI221D0 U2344 ( .A1(\entry[7][30] ), .A2(n2996), .B1(\entry[10][30] ), .B2(
        n2997), .C(n3140), .ZN(n3135) );
  AO22D0 U2345 ( .A1(\entry[6][30] ), .A2(n2999), .B1(\entry[5][30] ), .B2(
        n3000), .Z(n3140) );
  AOI221D0 U2346 ( .A1(\entry[14][30] ), .A2(n3001), .B1(\entry[9][30] ), .B2(
        n3002), .C(n3141), .ZN(n3134) );
  AO22D0 U2347 ( .A1(\entry[15][30] ), .A2(n3004), .B1(\entry[8][30] ), .B2(
        n3005), .Z(n3141) );
  ND4D0 U2348 ( .A1(n3142), .A2(n3143), .A3(n3144), .A4(n3145), .ZN(N10297) );
  AOI221D0 U2349 ( .A1(\entry[12][29] ), .A2(n2986), .B1(\entry[13][29] ), 
        .B2(n2987), .C(n3146), .ZN(n3145) );
  AO22D0 U2350 ( .A1(\entry[11][29] ), .A2(n2989), .B1(\entry[0][29] ), .B2(
        n2990), .Z(n3146) );
  AOI221D0 U2351 ( .A1(\entry[1][29] ), .A2(n2991), .B1(\entry[2][29] ), .B2(
        n2992), .C(n3147), .ZN(n3144) );
  AO22D0 U2352 ( .A1(\entry[4][29] ), .A2(n2994), .B1(\entry[3][29] ), .B2(
        n2995), .Z(n3147) );
  AOI221D0 U2353 ( .A1(\entry[7][29] ), .A2(n2996), .B1(\entry[10][29] ), .B2(
        n2997), .C(n3148), .ZN(n3143) );
  AO22D0 U2354 ( .A1(\entry[6][29] ), .A2(n2999), .B1(\entry[5][29] ), .B2(
        n3000), .Z(n3148) );
  AOI221D0 U2355 ( .A1(\entry[14][29] ), .A2(n3001), .B1(\entry[9][29] ), .B2(
        n3002), .C(n3149), .ZN(n3142) );
  AO22D0 U2356 ( .A1(\entry[15][29] ), .A2(n3004), .B1(\entry[8][29] ), .B2(
        n3005), .Z(n3149) );
  ND4D0 U2357 ( .A1(n3150), .A2(n3151), .A3(n3152), .A4(n3153), .ZN(N10296) );
  AOI221D0 U2358 ( .A1(\entry[12][28] ), .A2(n2986), .B1(\entry[13][28] ), 
        .B2(n2987), .C(n3154), .ZN(n3153) );
  AO22D0 U2359 ( .A1(\entry[11][28] ), .A2(n2989), .B1(\entry[0][28] ), .B2(
        n2990), .Z(n3154) );
  AOI221D0 U2360 ( .A1(\entry[1][28] ), .A2(n2991), .B1(\entry[2][28] ), .B2(
        n2992), .C(n3155), .ZN(n3152) );
  AO22D0 U2361 ( .A1(\entry[4][28] ), .A2(n2994), .B1(\entry[3][28] ), .B2(
        n2995), .Z(n3155) );
  AOI221D0 U2362 ( .A1(\entry[7][28] ), .A2(n2996), .B1(\entry[10][28] ), .B2(
        n2997), .C(n3156), .ZN(n3151) );
  AO22D0 U2363 ( .A1(\entry[6][28] ), .A2(n2999), .B1(\entry[5][28] ), .B2(
        n3000), .Z(n3156) );
  AOI221D0 U2364 ( .A1(\entry[14][28] ), .A2(n3001), .B1(\entry[9][28] ), .B2(
        n3002), .C(n3157), .ZN(n3150) );
  AO22D0 U2365 ( .A1(\entry[15][28] ), .A2(n3004), .B1(\entry[8][28] ), .B2(
        n3005), .Z(n3157) );
  ND4D0 U2366 ( .A1(n3158), .A2(n3159), .A3(n3160), .A4(n3161), .ZN(N10295) );
  AOI221D0 U2367 ( .A1(\entry[12][27] ), .A2(n2986), .B1(\entry[13][27] ), 
        .B2(n2987), .C(n3162), .ZN(n3161) );
  AO22D0 U2368 ( .A1(\entry[11][27] ), .A2(n2989), .B1(\entry[0][27] ), .B2(
        n2990), .Z(n3162) );
  AOI221D0 U2369 ( .A1(\entry[1][27] ), .A2(n2991), .B1(\entry[2][27] ), .B2(
        n2992), .C(n3163), .ZN(n3160) );
  AO22D0 U2370 ( .A1(\entry[4][27] ), .A2(n2994), .B1(\entry[3][27] ), .B2(
        n2995), .Z(n3163) );
  AOI221D0 U2371 ( .A1(\entry[7][27] ), .A2(n2996), .B1(\entry[10][27] ), .B2(
        n2997), .C(n3164), .ZN(n3159) );
  AO22D0 U2372 ( .A1(\entry[6][27] ), .A2(n2999), .B1(\entry[5][27] ), .B2(
        n3000), .Z(n3164) );
  AOI221D0 U2373 ( .A1(\entry[14][27] ), .A2(n3001), .B1(\entry[9][27] ), .B2(
        n3002), .C(n3165), .ZN(n3158) );
  AO22D0 U2374 ( .A1(\entry[15][27] ), .A2(n3004), .B1(\entry[8][27] ), .B2(
        n3005), .Z(n3165) );
  ND4D0 U2375 ( .A1(n3166), .A2(n3167), .A3(n3168), .A4(n3169), .ZN(N10294) );
  AOI221D0 U2376 ( .A1(\entry[12][26] ), .A2(n2986), .B1(\entry[13][26] ), 
        .B2(n2987), .C(n3170), .ZN(n3169) );
  AO22D0 U2377 ( .A1(\entry[11][26] ), .A2(n2989), .B1(\entry[0][26] ), .B2(
        n2990), .Z(n3170) );
  AOI221D0 U2378 ( .A1(\entry[1][26] ), .A2(n2991), .B1(\entry[2][26] ), .B2(
        n2992), .C(n3171), .ZN(n3168) );
  AO22D0 U2379 ( .A1(\entry[4][26] ), .A2(n2994), .B1(\entry[3][26] ), .B2(
        n2995), .Z(n3171) );
  AOI221D0 U2380 ( .A1(\entry[7][26] ), .A2(n2996), .B1(\entry[10][26] ), .B2(
        n2997), .C(n3172), .ZN(n3167) );
  AO22D0 U2381 ( .A1(\entry[6][26] ), .A2(n2999), .B1(\entry[5][26] ), .B2(
        n3000), .Z(n3172) );
  AOI221D0 U2382 ( .A1(\entry[14][26] ), .A2(n3001), .B1(\entry[9][26] ), .B2(
        n3002), .C(n3173), .ZN(n3166) );
  AO22D0 U2383 ( .A1(\entry[15][26] ), .A2(n3004), .B1(\entry[8][26] ), .B2(
        n3005), .Z(n3173) );
  ND4D0 U2384 ( .A1(n3174), .A2(n3175), .A3(n3176), .A4(n3177), .ZN(N10293) );
  AOI221D0 U2385 ( .A1(\entry[12][25] ), .A2(n2986), .B1(\entry[13][25] ), 
        .B2(n2987), .C(n3178), .ZN(n3177) );
  AO22D0 U2386 ( .A1(\entry[11][25] ), .A2(n2989), .B1(\entry[0][25] ), .B2(
        n2990), .Z(n3178) );
  AOI221D0 U2387 ( .A1(\entry[1][25] ), .A2(n2991), .B1(\entry[2][25] ), .B2(
        n2992), .C(n3179), .ZN(n3176) );
  AO22D0 U2388 ( .A1(\entry[4][25] ), .A2(n2994), .B1(\entry[3][25] ), .B2(
        n2995), .Z(n3179) );
  AOI221D0 U2389 ( .A1(\entry[7][25] ), .A2(n2996), .B1(\entry[10][25] ), .B2(
        n2997), .C(n3180), .ZN(n3175) );
  AO22D0 U2390 ( .A1(\entry[6][25] ), .A2(n2999), .B1(\entry[5][25] ), .B2(
        n3000), .Z(n3180) );
  AOI221D0 U2391 ( .A1(\entry[14][25] ), .A2(n3001), .B1(\entry[9][25] ), .B2(
        n3002), .C(n3181), .ZN(n3174) );
  AO22D0 U2392 ( .A1(\entry[15][25] ), .A2(n3004), .B1(\entry[8][25] ), .B2(
        n3005), .Z(n3181) );
  ND4D0 U2393 ( .A1(n3182), .A2(n3183), .A3(n3184), .A4(n3185), .ZN(N10292) );
  AOI221D0 U2394 ( .A1(\entry[12][24] ), .A2(n2986), .B1(\entry[13][24] ), 
        .B2(n2987), .C(n3186), .ZN(n3185) );
  AO22D0 U2395 ( .A1(\entry[11][24] ), .A2(n2989), .B1(\entry[0][24] ), .B2(
        n2990), .Z(n3186) );
  AOI221D0 U2396 ( .A1(\entry[1][24] ), .A2(n2991), .B1(\entry[2][24] ), .B2(
        n2992), .C(n3187), .ZN(n3184) );
  AO22D0 U2397 ( .A1(\entry[4][24] ), .A2(n2994), .B1(\entry[3][24] ), .B2(
        n2995), .Z(n3187) );
  AOI221D0 U2398 ( .A1(\entry[7][24] ), .A2(n2996), .B1(\entry[10][24] ), .B2(
        n2997), .C(n3188), .ZN(n3183) );
  AO22D0 U2399 ( .A1(\entry[6][24] ), .A2(n2999), .B1(\entry[5][24] ), .B2(
        n3000), .Z(n3188) );
  AOI221D0 U2400 ( .A1(\entry[14][24] ), .A2(n3001), .B1(\entry[9][24] ), .B2(
        n3002), .C(n3189), .ZN(n3182) );
  AO22D0 U2401 ( .A1(\entry[15][24] ), .A2(n3004), .B1(\entry[8][24] ), .B2(
        n3005), .Z(n3189) );
  ND4D0 U2402 ( .A1(n3190), .A2(n3191), .A3(n3192), .A4(n3193), .ZN(N10291) );
  AOI221D0 U2403 ( .A1(\entry[12][23] ), .A2(n2986), .B1(\entry[13][23] ), 
        .B2(n2987), .C(n3194), .ZN(n3193) );
  AO22D0 U2404 ( .A1(\entry[11][23] ), .A2(n2989), .B1(\entry[0][23] ), .B2(
        n2990), .Z(n3194) );
  AOI221D0 U2405 ( .A1(\entry[1][23] ), .A2(n2991), .B1(\entry[2][23] ), .B2(
        n2992), .C(n3195), .ZN(n3192) );
  AO22D0 U2406 ( .A1(\entry[4][23] ), .A2(n2994), .B1(\entry[3][23] ), .B2(
        n2995), .Z(n3195) );
  AOI221D0 U2407 ( .A1(\entry[7][23] ), .A2(n2996), .B1(\entry[10][23] ), .B2(
        n2997), .C(n3196), .ZN(n3191) );
  AO22D0 U2408 ( .A1(\entry[6][23] ), .A2(n2999), .B1(\entry[5][23] ), .B2(
        n3000), .Z(n3196) );
  AOI221D0 U2409 ( .A1(\entry[14][23] ), .A2(n3001), .B1(\entry[9][23] ), .B2(
        n3002), .C(n3197), .ZN(n3190) );
  AO22D0 U2410 ( .A1(\entry[15][23] ), .A2(n3004), .B1(\entry[8][23] ), .B2(
        n3005), .Z(n3197) );
  ND4D0 U2411 ( .A1(n3198), .A2(n3199), .A3(n3200), .A4(n3201), .ZN(N10290) );
  AOI221D0 U2412 ( .A1(\entry[12][22] ), .A2(n2986), .B1(\entry[13][22] ), 
        .B2(n2987), .C(n3202), .ZN(n3201) );
  AO22D0 U2413 ( .A1(\entry[11][22] ), .A2(n2989), .B1(\entry[0][22] ), .B2(
        n2990), .Z(n3202) );
  AOI221D0 U2414 ( .A1(\entry[1][22] ), .A2(n2991), .B1(\entry[2][22] ), .B2(
        n2992), .C(n3203), .ZN(n3200) );
  AO22D0 U2415 ( .A1(\entry[4][22] ), .A2(n2994), .B1(\entry[3][22] ), .B2(
        n2995), .Z(n3203) );
  AOI221D0 U2416 ( .A1(\entry[7][22] ), .A2(n2996), .B1(\entry[10][22] ), .B2(
        n2997), .C(n3204), .ZN(n3199) );
  AO22D0 U2417 ( .A1(\entry[6][22] ), .A2(n2999), .B1(\entry[5][22] ), .B2(
        n3000), .Z(n3204) );
  AOI221D0 U2418 ( .A1(\entry[14][22] ), .A2(n3001), .B1(\entry[9][22] ), .B2(
        n3002), .C(n3205), .ZN(n3198) );
  AO22D0 U2419 ( .A1(\entry[15][22] ), .A2(n3004), .B1(\entry[8][22] ), .B2(
        n3005), .Z(n3205) );
  ND4D0 U2420 ( .A1(n3206), .A2(n3207), .A3(n3208), .A4(n3209), .ZN(N10289) );
  AOI221D0 U2421 ( .A1(\entry[12][21] ), .A2(n2986), .B1(\entry[13][21] ), 
        .B2(n2987), .C(n3210), .ZN(n3209) );
  AO22D0 U2422 ( .A1(\entry[11][21] ), .A2(n2989), .B1(\entry[0][21] ), .B2(
        n2990), .Z(n3210) );
  AOI221D0 U2423 ( .A1(\entry[1][21] ), .A2(n2991), .B1(\entry[2][21] ), .B2(
        n2992), .C(n3211), .ZN(n3208) );
  AO22D0 U2424 ( .A1(\entry[4][21] ), .A2(n2994), .B1(\entry[3][21] ), .B2(
        n2995), .Z(n3211) );
  AOI221D0 U2425 ( .A1(\entry[7][21] ), .A2(n2996), .B1(\entry[10][21] ), .B2(
        n2997), .C(n3212), .ZN(n3207) );
  AO22D0 U2426 ( .A1(\entry[6][21] ), .A2(n2999), .B1(\entry[5][21] ), .B2(
        n3000), .Z(n3212) );
  AOI221D0 U2427 ( .A1(\entry[14][21] ), .A2(n3001), .B1(\entry[9][21] ), .B2(
        n3002), .C(n3213), .ZN(n3206) );
  AO22D0 U2428 ( .A1(\entry[15][21] ), .A2(n3004), .B1(\entry[8][21] ), .B2(
        n3005), .Z(n3213) );
  ND4D0 U2429 ( .A1(n3214), .A2(n3215), .A3(n3216), .A4(n3217), .ZN(N10288) );
  AOI221D0 U2430 ( .A1(\entry[12][20] ), .A2(n2986), .B1(\entry[13][20] ), 
        .B2(n2987), .C(n3218), .ZN(n3217) );
  AO22D0 U2431 ( .A1(\entry[11][20] ), .A2(n2989), .B1(\entry[0][20] ), .B2(
        n2990), .Z(n3218) );
  AOI221D0 U2432 ( .A1(\entry[1][20] ), .A2(n2991), .B1(\entry[2][20] ), .B2(
        n2992), .C(n3219), .ZN(n3216) );
  AO22D0 U2433 ( .A1(\entry[4][20] ), .A2(n2994), .B1(\entry[3][20] ), .B2(
        n2995), .Z(n3219) );
  AOI221D0 U2434 ( .A1(\entry[7][20] ), .A2(n2996), .B1(\entry[10][20] ), .B2(
        n2997), .C(n3220), .ZN(n3215) );
  AO22D0 U2435 ( .A1(\entry[6][20] ), .A2(n2999), .B1(\entry[5][20] ), .B2(
        n3000), .Z(n3220) );
  AOI221D0 U2436 ( .A1(\entry[14][20] ), .A2(n3001), .B1(\entry[9][20] ), .B2(
        n3002), .C(n3221), .ZN(n3214) );
  AO22D0 U2437 ( .A1(\entry[15][20] ), .A2(n3004), .B1(\entry[8][20] ), .B2(
        n3005), .Z(n3221) );
  ND4D0 U2438 ( .A1(n3222), .A2(n3223), .A3(n3224), .A4(n3225), .ZN(N10287) );
  AOI221D0 U2439 ( .A1(\entry[12][19] ), .A2(n2986), .B1(\entry[13][19] ), 
        .B2(n2987), .C(n3226), .ZN(n3225) );
  AO22D0 U2440 ( .A1(\entry[11][19] ), .A2(n2989), .B1(\entry[0][19] ), .B2(
        n2990), .Z(n3226) );
  AOI221D0 U2441 ( .A1(\entry[1][19] ), .A2(n2991), .B1(\entry[2][19] ), .B2(
        n2992), .C(n3227), .ZN(n3224) );
  AO22D0 U2442 ( .A1(\entry[4][19] ), .A2(n2994), .B1(\entry[3][19] ), .B2(
        n2995), .Z(n3227) );
  AOI221D0 U2443 ( .A1(\entry[7][19] ), .A2(n2996), .B1(\entry[10][19] ), .B2(
        n2997), .C(n3228), .ZN(n3223) );
  AO22D0 U2444 ( .A1(\entry[6][19] ), .A2(n2999), .B1(\entry[5][19] ), .B2(
        n3000), .Z(n3228) );
  AOI221D0 U2445 ( .A1(\entry[14][19] ), .A2(n3001), .B1(\entry[9][19] ), .B2(
        n3002), .C(n3229), .ZN(n3222) );
  AO22D0 U2446 ( .A1(\entry[15][19] ), .A2(n3004), .B1(\entry[8][19] ), .B2(
        n3005), .Z(n3229) );
  ND4D0 U2447 ( .A1(n3230), .A2(n3231), .A3(n3232), .A4(n3233), .ZN(N10286) );
  AOI221D0 U2448 ( .A1(\entry[12][18] ), .A2(n2986), .B1(\entry[13][18] ), 
        .B2(n2987), .C(n3234), .ZN(n3233) );
  AO22D0 U2449 ( .A1(\entry[11][18] ), .A2(n2989), .B1(\entry[0][18] ), .B2(
        n2990), .Z(n3234) );
  AOI221D0 U2450 ( .A1(\entry[1][18] ), .A2(n2991), .B1(\entry[2][18] ), .B2(
        n2992), .C(n3235), .ZN(n3232) );
  AO22D0 U2451 ( .A1(\entry[4][18] ), .A2(n2994), .B1(\entry[3][18] ), .B2(
        n2995), .Z(n3235) );
  AOI221D0 U2452 ( .A1(\entry[7][18] ), .A2(n2996), .B1(\entry[10][18] ), .B2(
        n2997), .C(n3236), .ZN(n3231) );
  AO22D0 U2453 ( .A1(\entry[6][18] ), .A2(n2999), .B1(\entry[5][18] ), .B2(
        n3000), .Z(n3236) );
  AOI221D0 U2454 ( .A1(\entry[14][18] ), .A2(n3001), .B1(\entry[9][18] ), .B2(
        n3002), .C(n3237), .ZN(n3230) );
  AO22D0 U2455 ( .A1(\entry[15][18] ), .A2(n3004), .B1(\entry[8][18] ), .B2(
        n3005), .Z(n3237) );
  ND4D0 U2456 ( .A1(n3238), .A2(n3239), .A3(n3240), .A4(n3241), .ZN(N10285) );
  AOI221D0 U2457 ( .A1(\entry[12][17] ), .A2(n2986), .B1(\entry[13][17] ), 
        .B2(n2987), .C(n3242), .ZN(n3241) );
  AO22D0 U2458 ( .A1(\entry[11][17] ), .A2(n2989), .B1(\entry[0][17] ), .B2(
        n2990), .Z(n3242) );
  CKND0 U2459 ( .I(n3246), .ZN(n3245) );
  AOI221D0 U2460 ( .A1(\entry[1][17] ), .A2(n2991), .B1(\entry[2][17] ), .B2(
        n2992), .C(n3247), .ZN(n3240) );
  AO22D0 U2461 ( .A1(\entry[4][17] ), .A2(n2994), .B1(\entry[3][17] ), .B2(
        n2995), .Z(n3247) );
  CKND0 U2462 ( .I(n3254), .ZN(n3253) );
  CKND0 U2463 ( .I(n3257), .ZN(n3256) );
  AOI221D0 U2464 ( .A1(\entry[7][17] ), .A2(n2996), .B1(\entry[10][17] ), .B2(
        n2997), .C(n3258), .ZN(n3239) );
  AO22D0 U2465 ( .A1(\entry[6][17] ), .A2(n2999), .B1(\entry[5][17] ), .B2(
        n3000), .Z(n3258) );
  AOI221D0 U2466 ( .A1(\entry[14][17] ), .A2(n3001), .B1(\entry[9][17] ), .B2(
        n3002), .C(n3265), .ZN(n3238) );
  AO22D0 U2467 ( .A1(\entry[15][17] ), .A2(n3004), .B1(\entry[8][17] ), .B2(
        n3005), .Z(n3265) );
  AN2D0 U2468 ( .A1(n3272), .A2(n3273), .Z(n3001) );
  OAI31D0 U2469 ( .A1(n3267), .A2(n3274), .A3(n3275), .B(n3243), .ZN(n3272) );
  ND4D0 U2470 ( .A1(n3276), .A2(n3277), .A3(n3278), .A4(n3279), .ZN(N10284) );
  AOI221D0 U2471 ( .A1(\entry[12][16] ), .A2(n2986), .B1(\entry[13][16] ), 
        .B2(n2987), .C(n3280), .ZN(n3279) );
  AO22D0 U2472 ( .A1(\entry[11][16] ), .A2(n2989), .B1(n3281), .B2(n3282), .Z(
        n3280) );
  OAI22D0 U2473 ( .A1(n3271), .A2(n3283), .B1(n3284), .B2(n3285), .ZN(n3282)
         );
  AOI32D0 U2474 ( .A1(\entry[14][16] ), .A2(n3286), .A3(n3287), .B1(
        \entry[8][16] ), .B2(n3288), .ZN(n3284) );
  INR2D0 U2475 ( .A1(n3273), .B1(n3274), .ZN(n3287) );
  CKND0 U2476 ( .I(n3275), .ZN(n3286) );
  OA21D0 U2477 ( .A1(n3291), .A2(n3292), .B(n3293), .Z(n2989) );
  NR2D0 U2478 ( .A1(n3243), .A2(n3294), .ZN(n3291) );
  AN2D0 U2479 ( .A1(n3295), .A2(n3274), .Z(n2987) );
  OAI22D0 U2480 ( .A1(n3273), .A2(n3243), .B1(n3275), .B2(n3267), .ZN(n3295)
         );
  AN2D0 U2481 ( .A1(n3296), .A2(n3297), .Z(n2986) );
  OAI32D0 U2482 ( .A1(n3243), .A2(n3274), .A3(n3273), .B1(n3293), .B2(n3298), 
        .ZN(n3296) );
  CKND0 U2483 ( .I(n3292), .ZN(n3298) );
  NR4D0 U2484 ( .A1(n3267), .A2(n3288), .A3(n3289), .A4(n3299), .ZN(n3292) );
  AOI221D0 U2485 ( .A1(\entry[10][16] ), .A2(n2997), .B1(\entry[1][16] ), .B2(
        n3257), .C(n3300), .ZN(n3278) );
  OAI22D0 U2486 ( .A1(n3260), .A2(n3301), .B1(n3249), .B2(n3302), .ZN(n3300)
         );
  ND4D0 U2487 ( .A1(n3281), .A2(n3303), .A3(n3304), .A4(n3305), .ZN(n3249) );
  IND3D0 U2488 ( .A1(n3306), .B1(n3307), .B2(n3308), .ZN(n3260) );
  NR2D0 U2489 ( .A1(n3270), .A2(n3304), .ZN(n3257) );
  CKND0 U2490 ( .I(n3309), .ZN(n3304) );
  AN2D0 U2491 ( .A1(n3310), .A2(n3299), .Z(n2997) );
  OAI33D0 U2492 ( .A1(n3294), .A2(n3293), .A3(n3243), .B1(n3267), .B2(n3289), 
        .B3(n3288), .ZN(n3310) );
  CKND2D0 U2493 ( .A1(n3281), .A2(n3290), .ZN(n3267) );
  CKND0 U2494 ( .I(n3311), .ZN(n3294) );
  AOI221D0 U2495 ( .A1(n3246), .A2(\entry[0][16] ), .B1(n3312), .B2(
        \entry[4][16] ), .C(n3313), .ZN(n3277) );
  OAI22D0 U2496 ( .A1(n3314), .A2(n3264), .B1(n3315), .B2(n3243), .ZN(n3313)
         );
  CKND2D0 U2497 ( .A1(val[15]), .A2(n3316), .ZN(n3243) );
  NR4D0 U2498 ( .A1(n3317), .A2(n3318), .A3(n3319), .A4(n3320), .ZN(n3315) );
  MOAI22D0 U2499 ( .A1(n3244), .A2(n3321), .B1(n3273), .B2(\entry[14][16] ), 
        .ZN(n3320) );
  CKND0 U2500 ( .I(\entry[0][16] ), .ZN(n3321) );
  OAI222D0 U2501 ( .A1(n3259), .A2(n3301), .B1(n3261), .B2(n3322), .C1(n3269), 
        .C2(n3283), .ZN(n3319) );
  CKND0 U2502 ( .I(\entry[9][16] ), .ZN(n3283) );
  IIND4D0 U2503 ( .A1(n3293), .A2(n3299), .B1(n3311), .B2(n3289), .ZN(n3269)
         );
  CKND0 U2504 ( .I(\entry[6][16] ), .ZN(n3322) );
  IND3D0 U2505 ( .A1(n3323), .B1(n3324), .B2(n3325), .ZN(n3261) );
  CKND0 U2506 ( .I(\entry[5][16] ), .ZN(n3301) );
  ND3D0 U2507 ( .A1(n3326), .A2(n3307), .A3(n3325), .ZN(n3259) );
  OAI222D0 U2508 ( .A1(n3255), .A2(n3327), .B1(n3250), .B2(n3328), .C1(n3248), 
        .C2(n3302), .ZN(n3318) );
  CKND0 U2509 ( .I(\entry[3][16] ), .ZN(n3302) );
  ND3D0 U2510 ( .A1(n3325), .A2(n3305), .A3(n3329), .ZN(n3248) );
  CKND0 U2511 ( .I(\entry[4][16] ), .ZN(n3328) );
  IND4D0 U2512 ( .A1(n3307), .B1(n3325), .B2(n3326), .B3(n3306), .ZN(n3250) );
  CKND0 U2513 ( .I(\entry[1][16] ), .ZN(n3327) );
  ND3D0 U2514 ( .A1(n3303), .A2(n3309), .A3(n3330), .ZN(n3255) );
  OAI222D0 U2515 ( .A1(n3263), .A2(n3314), .B1(n3268), .B2(n3331), .C1(n3252), 
        .C2(n3332), .ZN(n3317) );
  CKND0 U2516 ( .I(\entry[2][16] ), .ZN(n3332) );
  CKND2D0 U2517 ( .A1(n3330), .A2(n3333), .ZN(n3252) );
  CKND0 U2518 ( .I(n3334), .ZN(n3330) );
  IND3D0 U2519 ( .A1(n3305), .B1(n3325), .B2(n3329), .ZN(n3334) );
  INR3D0 U2520 ( .A1(n3326), .B1(n3307), .B2(n3306), .ZN(n3329) );
  CKND0 U2521 ( .I(\entry[8][16] ), .ZN(n3331) );
  ND3D0 U2522 ( .A1(n3335), .A2(n3288), .A3(n3311), .ZN(n3268) );
  NR3D0 U2523 ( .A1(n3274), .A2(n3297), .A3(n3273), .ZN(n3311) );
  CKND2D0 U2524 ( .A1(n3325), .A2(n3323), .ZN(n3263) );
  IND4D0 U2525 ( .A1(n3324), .B1(n3281), .B2(n3336), .B3(n3323), .ZN(n3264) );
  CKND0 U2526 ( .I(\entry[7][16] ), .ZN(n3314) );
  CKND0 U2527 ( .I(n3251), .ZN(n3312) );
  CKND2D0 U2528 ( .A1(n3308), .A2(n3306), .ZN(n3251) );
  NR4D0 U2529 ( .A1(n3270), .A2(n3305), .A3(n3333), .A4(n3309), .ZN(n3308) );
  AOI21D0 U2530 ( .A1(n3343), .A2(n3342), .B(val[15]), .ZN(n3246) );
  AOI222D0 U2531 ( .A1(n3337), .A2(\entry[6][16] ), .B1(\entry[15][16] ), .B2(
        n3004), .C1(n3254), .C2(\entry[2][16] ), .ZN(n3276) );
  NR3D0 U2532 ( .A1(n3309), .A2(n3303), .A3(n3270), .ZN(n3254) );
  CKND0 U2533 ( .I(n3333), .ZN(n3303) );
  AN2D0 U2534 ( .A1(n3340), .A2(n3341), .Z(n3316) );
  CKND2D0 U2535 ( .A1(n3290), .A2(n3325), .ZN(n3244) );
  NR3D0 U2536 ( .A1(n3273), .A2(n3274), .A3(n3275), .ZN(n3325) );
  IND3D0 U2537 ( .A1(n3297), .B1(n3335), .B2(n3266), .ZN(n3275) );
  CKND0 U2538 ( .I(n3288), .ZN(n3266) );
  CKND2D0 U2539 ( .A1(n2189), .A2(n2190), .ZN(n3288) );
  NR3D0 U2540 ( .A1(n3299), .A2(n3293), .A3(n3289), .ZN(n3335) );
  CKND2D0 U2541 ( .A1(n2191), .A2(n2192), .ZN(n3289) );
  CKND2D0 U2542 ( .A1(n2187), .A2(n2188), .ZN(n3293) );
  CKND2D0 U2543 ( .A1(n2193), .A2(n2194), .ZN(n3299) );
  CKND2D0 U2544 ( .A1(n2185), .A2(n2186), .ZN(n3297) );
  CKND2D0 U2545 ( .A1(n2184), .A2(n2183), .ZN(n3274) );
  CKND2D0 U2546 ( .A1(n2181), .A2(n2182), .ZN(n3273) );
  CKND0 U2547 ( .I(n3285), .ZN(n3290) );
  CKND2D0 U2548 ( .A1(n3336), .A2(n3326), .ZN(n3285) );
  NR2D0 U2549 ( .A1(n3324), .A2(n3323), .ZN(n3326) );
  CKND2D0 U2550 ( .A1(n2195), .A2(n2196), .ZN(n3323) );
  CKND0 U2551 ( .I(n3262), .ZN(n3337) );
  ND3D0 U2552 ( .A1(n3336), .A2(n3324), .A3(n3281), .ZN(n3262) );
  CKND0 U2553 ( .I(n3270), .ZN(n3281) );
  ND3D0 U2554 ( .A1(n3343), .A2(n3338), .A3(n3342), .ZN(n3270) );
  CKND0 U2555 ( .I(val[15]), .ZN(n3338) );
  CKND2D0 U2556 ( .A1(n2197), .A2(n2198), .ZN(n3324) );
  INR4D0 U2557 ( .A1(n3339), .B1(n3309), .B2(n3306), .B3(n3333), .ZN(n3336) );
  CKND2D0 U2558 ( .A1(n2205), .A2(n2206), .ZN(n3333) );
  CKND2D0 U2559 ( .A1(n2201), .A2(n2202), .ZN(n3306) );
  CKND2D0 U2560 ( .A1(n2203), .A2(n2204), .ZN(n3309) );
  NR2D0 U2561 ( .A1(n3305), .A2(n3307), .ZN(n3339) );
  CKND2D0 U2562 ( .A1(n2199), .A2(n2200), .ZN(n3307) );
  CKND2D0 U2563 ( .A1(n2207), .A2(n2208), .ZN(n3305) );
endmodule

